// mem_cp.v
// to be included from the top module at the compile

initial
begin
mem_cp['o0000]='o0000;
mem_cp['o0001]='o0000;
mem_cp['o0002]='o0000;
mem_cp['o0003]='o0000;
mem_cp['o0004]='o0000;
mem_cp['o0005]='o0000;
mem_cp['o0006]='o0000;
mem_cp['o0007]='o0000;
mem_cp['o0010]='o0000;
mem_cp['o0011]='o0000;
mem_cp['o0012]='o0000;
mem_cp['o0013]='o0000;
mem_cp['o0014]='o0000;
mem_cp['o0015]='o0000;
mem_cp['o0016]='o0000;
mem_cp['o0017]='o0000;
mem_cp['o0020]='o0000;
mem_cp['o0021]='o0000;
mem_cp['o0022]='o0000;
mem_cp['o0023]='o0000;
mem_cp['o0024]='o0000;
mem_cp['o0025]='o0000;
mem_cp['o0026]='o0000;
mem_cp['o0027]='o0000;
mem_cp['o0030]='o0000;
mem_cp['o0031]='o0000;
mem_cp['o0032]='o0000;
mem_cp['o0033]='o0000;
mem_cp['o0034]='o0000;
mem_cp['o0035]='o0000;
mem_cp['o0036]='o0000;
mem_cp['o0037]='o0000;
mem_cp['o0040]='o0000;
mem_cp['o0041]='o0000;
mem_cp['o0042]='o0000;
mem_cp['o0043]='o0000;
mem_cp['o0044]='o0000;
mem_cp['o0045]='o0000;
mem_cp['o0046]='o0000;
mem_cp['o0047]='o0000;
mem_cp['o0050]='o0000;
mem_cp['o0051]='o0000;
mem_cp['o0052]='o0000;
mem_cp['o0053]='o0000;
mem_cp['o0054]='o0000;
mem_cp['o0055]='o0000;
mem_cp['o0056]='o0000;
mem_cp['o0057]='o0000;
mem_cp['o0060]='o0000;
mem_cp['o0061]='o0000;
mem_cp['o0062]='o0000;
mem_cp['o0063]='o0000;
mem_cp['o0064]='o0000;
mem_cp['o0065]='o0000;
mem_cp['o0066]='o0000;
mem_cp['o0067]='o0000;
mem_cp['o0070]='o0000;
mem_cp['o0071]='o0000;
mem_cp['o0072]='o0000;
mem_cp['o0073]='o0000;
mem_cp['o0074]='o0000;
mem_cp['o0075]='o0000;
mem_cp['o0076]='o0000;
mem_cp['o0077]='o0000;
mem_cp['o0100]='o5000;
mem_cp['o0101]='o5046;
mem_cp['o0102]='o7423;
mem_cp['o0103]='o7200;
mem_cp['o0104]='o7405;
mem_cp['o0105]='o7414;
mem_cp['o0106]='o0000;
mem_cp['o0107]='o5111;
mem_cp['o0110]='o7000;
mem_cp['o0111]='o7014;
mem_cp['o0112]='o7032;
mem_cp['o0113]='o6646;
mem_cp['o0114]='o6620;
mem_cp['o0115]='o6634;
mem_cp['o0116]='o0000;
mem_cp['o0117]='o0000;
mem_cp['o0120]='o0000;
mem_cp['o0121]='o0000;
mem_cp['o0122]='o0000;
mem_cp['o0123]='o0000;
mem_cp['o0124]='o0000;
mem_cp['o0125]='o0000;
mem_cp['o0126]='o0000;
mem_cp['o0127]='o0000;
mem_cp['o0130]='o0000;
mem_cp['o0131]='o0000;
mem_cp['o0132]='o0000;
mem_cp['o0133]='o0000;
mem_cp['o0134]='o0000;
mem_cp['o0135]='o0000;
mem_cp['o0136]='o0000;
mem_cp['o0137]='o0000;
mem_cp['o0140]='o0000;
mem_cp['o0141]='o0000;
mem_cp['o0142]='o0000;
mem_cp['o0143]='o0000;
mem_cp['o0144]='o0000;
mem_cp['o0145]='o0000;
mem_cp['o0146]='o0000;
mem_cp['o0147]='o0000;
mem_cp['o0150]='o0000;
mem_cp['o0151]='o0000;
mem_cp['o0152]='o1417;
mem_cp['o0153]='o7200;
mem_cp['o0154]='o1017;
mem_cp['o0155]='o1173;
mem_cp['o0156]='o3157;
mem_cp['o0157]='o7000;
mem_cp['o0160]='o5551;
mem_cp['o0161]='o0000;
mem_cp['o0162]='o7421;
mem_cp['o0163]='o1417;
mem_cp['o0164]='o7200;
mem_cp['o0165]='o1017;
mem_cp['o0166]='o1174;
mem_cp['o0167]='o3171;
mem_cp['o0170]='o7501;
mem_cp['o0171]='o7000;
mem_cp['o0172]='o5561;
mem_cp['o0173]='o1000;
mem_cp['o0174]='o3000;
mem_cp['o0175]='o0000;
mem_cp['o0176]='o0000;
mem_cp['o0177]='o0000;
mem_cp['o0200]='o0000;
mem_cp['o0201]='o0000;
mem_cp['o0202]='o0000;
mem_cp['o0203]='o0000;
mem_cp['o0204]='o0000;
mem_cp['o0205]='o0000;
mem_cp['o0206]='o0000;
mem_cp['o0207]='o0000;
mem_cp['o0210]='o0000;
mem_cp['o0211]='o0000;
mem_cp['o0212]='o0000;
mem_cp['o0213]='o0000;
mem_cp['o0214]='o0000;
mem_cp['o0215]='o0000;
mem_cp['o0216]='o0000;
mem_cp['o0217]='o0000;
mem_cp['o0220]='o0000;
mem_cp['o0221]='o0000;
mem_cp['o0222]='o0000;
mem_cp['o0223]='o0000;
mem_cp['o0224]='o0000;
mem_cp['o0225]='o0000;
mem_cp['o0226]='o0000;
mem_cp['o0227]='o0000;
mem_cp['o0230]='o0000;
mem_cp['o0231]='o0000;
mem_cp['o0232]='o0000;
mem_cp['o0233]='o0000;
mem_cp['o0234]='o0000;
mem_cp['o0235]='o0000;
mem_cp['o0236]='o0000;
mem_cp['o0237]='o0000;
mem_cp['o0240]='o0000;
mem_cp['o0241]='o0000;
mem_cp['o0242]='o0000;
mem_cp['o0243]='o0000;
mem_cp['o0244]='o0000;
mem_cp['o0245]='o0000;
mem_cp['o0246]='o0000;
mem_cp['o0247]='o0000;
mem_cp['o0250]='o0000;
mem_cp['o0251]='o0000;
mem_cp['o0252]='o0000;
mem_cp['o0253]='o0000;
mem_cp['o0254]='o0000;
mem_cp['o0255]='o0000;
mem_cp['o0256]='o0000;
mem_cp['o0257]='o0000;
mem_cp['o0260]='o0000;
mem_cp['o0261]='o0000;
mem_cp['o0262]='o0000;
mem_cp['o0263]='o0000;
mem_cp['o0264]='o0000;
mem_cp['o0265]='o0000;
mem_cp['o0266]='o0000;
mem_cp['o0267]='o0000;
mem_cp['o0270]='o0000;
mem_cp['o0271]='o0000;
mem_cp['o0272]='o0000;
mem_cp['o0273]='o0000;
mem_cp['o0274]='o0000;
mem_cp['o0275]='o0000;
mem_cp['o0276]='o0000;
mem_cp['o0277]='o0000;
mem_cp['o0300]='o0000;
mem_cp['o0301]='o0000;
mem_cp['o0302]='o0000;
mem_cp['o0303]='o0000;
mem_cp['o0304]='o0000;
mem_cp['o0305]='o0000;
mem_cp['o0306]='o0000;
mem_cp['o0307]='o0000;
mem_cp['o0310]='o0000;
mem_cp['o0311]='o0000;
mem_cp['o0312]='o0000;
mem_cp['o0313]='o0000;
mem_cp['o0314]='o0000;
mem_cp['o0315]='o0000;
mem_cp['o0316]='o0000;
mem_cp['o0317]='o0000;
mem_cp['o0320]='o0000;
mem_cp['o0321]='o0000;
mem_cp['o0322]='o0000;
mem_cp['o0323]='o0000;
mem_cp['o0324]='o0000;
mem_cp['o0325]='o0000;
mem_cp['o0326]='o0000;
mem_cp['o0327]='o0000;
mem_cp['o0330]='o0000;
mem_cp['o0331]='o0000;
mem_cp['o0332]='o0000;
mem_cp['o0333]='o0000;
mem_cp['o0334]='o0000;
mem_cp['o0335]='o0000;
mem_cp['o0336]='o0000;
mem_cp['o0337]='o0000;
mem_cp['o0340]='o0000;
mem_cp['o0341]='o0000;
mem_cp['o0342]='o0000;
mem_cp['o0343]='o0000;
mem_cp['o0344]='o0000;
mem_cp['o0345]='o0000;
mem_cp['o0346]='o0000;
mem_cp['o0347]='o0000;
mem_cp['o0350]='o0000;
mem_cp['o0351]='o0000;
mem_cp['o0352]='o0000;
mem_cp['o0353]='o0000;
mem_cp['o0354]='o0000;
mem_cp['o0355]='o0000;
mem_cp['o0356]='o0000;
mem_cp['o0357]='o0000;
mem_cp['o0360]='o0000;
mem_cp['o0361]='o0000;
mem_cp['o0362]='o0000;
mem_cp['o0363]='o0000;
mem_cp['o0364]='o0000;
mem_cp['o0365]='o0000;
mem_cp['o0366]='o0000;
mem_cp['o0367]='o0000;
mem_cp['o0370]='o0000;
mem_cp['o0371]='o0000;
mem_cp['o0372]='o0000;
mem_cp['o0373]='o0000;
mem_cp['o0374]='o0000;
mem_cp['o0375]='o0000;
mem_cp['o0376]='o0000;
mem_cp['o0377]='o0000;
mem_cp['o0400]='o0000;
mem_cp['o0401]='o0000;
mem_cp['o0402]='o0000;
mem_cp['o0403]='o0000;
mem_cp['o0404]='o0000;
mem_cp['o0405]='o0000;
mem_cp['o0406]='o0000;
mem_cp['o0407]='o0000;
mem_cp['o0410]='o0000;
mem_cp['o0411]='o0000;
mem_cp['o0412]='o0000;
mem_cp['o0413]='o0000;
mem_cp['o0414]='o0000;
mem_cp['o0415]='o0000;
mem_cp['o0416]='o0000;
mem_cp['o0417]='o0000;
mem_cp['o0420]='o0000;
mem_cp['o0421]='o0000;
mem_cp['o0422]='o0000;
mem_cp['o0423]='o0000;
mem_cp['o0424]='o0000;
mem_cp['o0425]='o0000;
mem_cp['o0426]='o0000;
mem_cp['o0427]='o0000;
mem_cp['o0430]='o0000;
mem_cp['o0431]='o0000;
mem_cp['o0432]='o0000;
mem_cp['o0433]='o0000;
mem_cp['o0434]='o0000;
mem_cp['o0435]='o0000;
mem_cp['o0436]='o0000;
mem_cp['o0437]='o0000;
mem_cp['o0440]='o0000;
mem_cp['o0441]='o0000;
mem_cp['o0442]='o0000;
mem_cp['o0443]='o0000;
mem_cp['o0444]='o0000;
mem_cp['o0445]='o0000;
mem_cp['o0446]='o0000;
mem_cp['o0447]='o0000;
mem_cp['o0450]='o0000;
mem_cp['o0451]='o0000;
mem_cp['o0452]='o0000;
mem_cp['o0453]='o0000;
mem_cp['o0454]='o0000;
mem_cp['o0455]='o0000;
mem_cp['o0456]='o0000;
mem_cp['o0457]='o0000;
mem_cp['o0460]='o0000;
mem_cp['o0461]='o0000;
mem_cp['o0462]='o0000;
mem_cp['o0463]='o0000;
mem_cp['o0464]='o0000;
mem_cp['o0465]='o0000;
mem_cp['o0466]='o0000;
mem_cp['o0467]='o0000;
mem_cp['o0470]='o0000;
mem_cp['o0471]='o0000;
mem_cp['o0472]='o0000;
mem_cp['o0473]='o0000;
mem_cp['o0474]='o0000;
mem_cp['o0475]='o0000;
mem_cp['o0476]='o0000;
mem_cp['o0477]='o0000;
mem_cp['o0500]='o0000;
mem_cp['o0501]='o0000;
mem_cp['o0502]='o0000;
mem_cp['o0503]='o0000;
mem_cp['o0504]='o0000;
mem_cp['o0505]='o0000;
mem_cp['o0506]='o0000;
mem_cp['o0507]='o0000;
mem_cp['o0510]='o0000;
mem_cp['o0511]='o0000;
mem_cp['o0512]='o0000;
mem_cp['o0513]='o0000;
mem_cp['o0514]='o0000;
mem_cp['o0515]='o0000;
mem_cp['o0516]='o0000;
mem_cp['o0517]='o0000;
mem_cp['o0520]='o0000;
mem_cp['o0521]='o0000;
mem_cp['o0522]='o0000;
mem_cp['o0523]='o0000;
mem_cp['o0524]='o0000;
mem_cp['o0525]='o0000;
mem_cp['o0526]='o0000;
mem_cp['o0527]='o0000;
mem_cp['o0530]='o0000;
mem_cp['o0531]='o0000;
mem_cp['o0532]='o0000;
mem_cp['o0533]='o0000;
mem_cp['o0534]='o0000;
mem_cp['o0535]='o0000;
mem_cp['o0536]='o0000;
mem_cp['o0537]='o0000;
mem_cp['o0540]='o0000;
mem_cp['o0541]='o0000;
mem_cp['o0542]='o0000;
mem_cp['o0543]='o0000;
mem_cp['o0544]='o0000;
mem_cp['o0545]='o0000;
mem_cp['o0546]='o0000;
mem_cp['o0547]='o0000;
mem_cp['o0550]='o0000;
mem_cp['o0551]='o0000;
mem_cp['o0552]='o0000;
mem_cp['o0553]='o0000;
mem_cp['o0554]='o0000;
mem_cp['o0555]='o0000;
mem_cp['o0556]='o0000;
mem_cp['o0557]='o0000;
mem_cp['o0560]='o0000;
mem_cp['o0561]='o0000;
mem_cp['o0562]='o0000;
mem_cp['o0563]='o0000;
mem_cp['o0564]='o0000;
mem_cp['o0565]='o0000;
mem_cp['o0566]='o0000;
mem_cp['o0567]='o0000;
mem_cp['o0570]='o0000;
mem_cp['o0571]='o0000;
mem_cp['o0572]='o0000;
mem_cp['o0573]='o0000;
mem_cp['o0574]='o0000;
mem_cp['o0575]='o0000;
mem_cp['o0576]='o0000;
mem_cp['o0577]='o0000;
mem_cp['o0600]='o0000;
mem_cp['o0601]='o0000;
mem_cp['o0602]='o0000;
mem_cp['o0603]='o0000;
mem_cp['o0604]='o0000;
mem_cp['o0605]='o0000;
mem_cp['o0606]='o0000;
mem_cp['o0607]='o0000;
mem_cp['o0610]='o0000;
mem_cp['o0611]='o0000;
mem_cp['o0612]='o0000;
mem_cp['o0613]='o0000;
mem_cp['o0614]='o0000;
mem_cp['o0615]='o0000;
mem_cp['o0616]='o0000;
mem_cp['o0617]='o0000;
mem_cp['o0620]='o0000;
mem_cp['o0621]='o0000;
mem_cp['o0622]='o0000;
mem_cp['o0623]='o0000;
mem_cp['o0624]='o0000;
mem_cp['o0625]='o0000;
mem_cp['o0626]='o0000;
mem_cp['o0627]='o0000;
mem_cp['o0630]='o0000;
mem_cp['o0631]='o0000;
mem_cp['o0632]='o0000;
mem_cp['o0633]='o0000;
mem_cp['o0634]='o0000;
mem_cp['o0635]='o0000;
mem_cp['o0636]='o0000;
mem_cp['o0637]='o0000;
mem_cp['o0640]='o0000;
mem_cp['o0641]='o0000;
mem_cp['o0642]='o0000;
mem_cp['o0643]='o0000;
mem_cp['o0644]='o0000;
mem_cp['o0645]='o0000;
mem_cp['o0646]='o0000;
mem_cp['o0647]='o0000;
mem_cp['o0650]='o0000;
mem_cp['o0651]='o0000;
mem_cp['o0652]='o0000;
mem_cp['o0653]='o0000;
mem_cp['o0654]='o0000;
mem_cp['o0655]='o0000;
mem_cp['o0656]='o0000;
mem_cp['o0657]='o0000;
mem_cp['o0660]='o0000;
mem_cp['o0661]='o0000;
mem_cp['o0662]='o0000;
mem_cp['o0663]='o0000;
mem_cp['o0664]='o0000;
mem_cp['o0665]='o0000;
mem_cp['o0666]='o0000;
mem_cp['o0667]='o0000;
mem_cp['o0670]='o0000;
mem_cp['o0671]='o0000;
mem_cp['o0672]='o0000;
mem_cp['o0673]='o0000;
mem_cp['o0674]='o0000;
mem_cp['o0675]='o0000;
mem_cp['o0676]='o0000;
mem_cp['o0677]='o0000;
mem_cp['o0700]='o0000;
mem_cp['o0701]='o0000;
mem_cp['o0702]='o0000;
mem_cp['o0703]='o0000;
mem_cp['o0704]='o0000;
mem_cp['o0705]='o0000;
mem_cp['o0706]='o0000;
mem_cp['o0707]='o0000;
mem_cp['o0710]='o0000;
mem_cp['o0711]='o0000;
mem_cp['o0712]='o0000;
mem_cp['o0713]='o0000;
mem_cp['o0714]='o0000;
mem_cp['o0715]='o0000;
mem_cp['o0716]='o0000;
mem_cp['o0717]='o0000;
mem_cp['o0720]='o0000;
mem_cp['o0721]='o0000;
mem_cp['o0722]='o0000;
mem_cp['o0723]='o0000;
mem_cp['o0724]='o0000;
mem_cp['o0725]='o0000;
mem_cp['o0726]='o0000;
mem_cp['o0727]='o0000;
mem_cp['o0730]='o0000;
mem_cp['o0731]='o0000;
mem_cp['o0732]='o0000;
mem_cp['o0733]='o0000;
mem_cp['o0734]='o0000;
mem_cp['o0735]='o0000;
mem_cp['o0736]='o0000;
mem_cp['o0737]='o0000;
mem_cp['o0740]='o0000;
mem_cp['o0741]='o0000;
mem_cp['o0742]='o0000;
mem_cp['o0743]='o0000;
mem_cp['o0744]='o0000;
mem_cp['o0745]='o0000;
mem_cp['o0746]='o0000;
mem_cp['o0747]='o0000;
mem_cp['o0750]='o0000;
mem_cp['o0751]='o0000;
mem_cp['o0752]='o0000;
mem_cp['o0753]='o0000;
mem_cp['o0754]='o0000;
mem_cp['o0755]='o0000;
mem_cp['o0756]='o0000;
mem_cp['o0757]='o0000;
mem_cp['o0760]='o0000;
mem_cp['o0761]='o0000;
mem_cp['o0762]='o0000;
mem_cp['o0763]='o0000;
mem_cp['o0764]='o0000;
mem_cp['o0765]='o0000;
mem_cp['o0766]='o0000;
mem_cp['o0767]='o0000;
mem_cp['o0770]='o0000;
mem_cp['o0771]='o0000;
mem_cp['o0772]='o0000;
mem_cp['o0773]='o0000;
mem_cp['o0774]='o0000;
mem_cp['o0775]='o0000;
mem_cp['o0776]='o0000;
mem_cp['o0777]='o0000;
mem_cp['o1000]='o0000;
mem_cp['o1001]='o0000;
mem_cp['o1002]='o0000;
mem_cp['o1003]='o0000;
mem_cp['o1004]='o0000;
mem_cp['o1005]='o0000;
mem_cp['o1006]='o0000;
mem_cp['o1007]='o0000;
mem_cp['o1010]='o0000;
mem_cp['o1011]='o0000;
mem_cp['o1012]='o0000;
mem_cp['o1013]='o0000;
mem_cp['o1014]='o0000;
mem_cp['o1015]='o0000;
mem_cp['o1016]='o0000;
mem_cp['o1017]='o0000;
mem_cp['o1020]='o0000;
mem_cp['o1021]='o0000;
mem_cp['o1022]='o0000;
mem_cp['o1023]='o0000;
mem_cp['o1024]='o0000;
mem_cp['o1025]='o0000;
mem_cp['o1026]='o0000;
mem_cp['o1027]='o0000;
mem_cp['o1030]='o0000;
mem_cp['o1031]='o0000;
mem_cp['o1032]='o0000;
mem_cp['o1033]='o0000;
mem_cp['o1034]='o0000;
mem_cp['o1035]='o0000;
mem_cp['o1036]='o0000;
mem_cp['o1037]='o0000;
mem_cp['o1040]='o0000;
mem_cp['o1041]='o0000;
mem_cp['o1042]='o0000;
mem_cp['o1043]='o0000;
mem_cp['o1044]='o0000;
mem_cp['o1045]='o0000;
mem_cp['o1046]='o0000;
mem_cp['o1047]='o0000;
mem_cp['o1050]='o0000;
mem_cp['o1051]='o0000;
mem_cp['o1052]='o0000;
mem_cp['o1053]='o0000;
mem_cp['o1054]='o0000;
mem_cp['o1055]='o0000;
mem_cp['o1056]='o0000;
mem_cp['o1057]='o0000;
mem_cp['o1060]='o0000;
mem_cp['o1061]='o0000;
mem_cp['o1062]='o0000;
mem_cp['o1063]='o0000;
mem_cp['o1064]='o0000;
mem_cp['o1065]='o0000;
mem_cp['o1066]='o0000;
mem_cp['o1067]='o0000;
mem_cp['o1070]='o0000;
mem_cp['o1071]='o0000;
mem_cp['o1072]='o0000;
mem_cp['o1073]='o0000;
mem_cp['o1074]='o0000;
mem_cp['o1075]='o0000;
mem_cp['o1076]='o0000;
mem_cp['o1077]='o0000;
mem_cp['o1100]='o0000;
mem_cp['o1101]='o0000;
mem_cp['o1102]='o0000;
mem_cp['o1103]='o0000;
mem_cp['o1104]='o0000;
mem_cp['o1105]='o0000;
mem_cp['o1106]='o0000;
mem_cp['o1107]='o0000;
mem_cp['o1110]='o0000;
mem_cp['o1111]='o0000;
mem_cp['o1112]='o0000;
mem_cp['o1113]='o0000;
mem_cp['o1114]='o0000;
mem_cp['o1115]='o0000;
mem_cp['o1116]='o0000;
mem_cp['o1117]='o0000;
mem_cp['o1120]='o0000;
mem_cp['o1121]='o0000;
mem_cp['o1122]='o0000;
mem_cp['o1123]='o0000;
mem_cp['o1124]='o0000;
mem_cp['o1125]='o0000;
mem_cp['o1126]='o0000;
mem_cp['o1127]='o0000;
mem_cp['o1130]='o0000;
mem_cp['o1131]='o0000;
mem_cp['o1132]='o0000;
mem_cp['o1133]='o0000;
mem_cp['o1134]='o0000;
mem_cp['o1135]='o0000;
mem_cp['o1136]='o0000;
mem_cp['o1137]='o0000;
mem_cp['o1140]='o0000;
mem_cp['o1141]='o0000;
mem_cp['o1142]='o0000;
mem_cp['o1143]='o0000;
mem_cp['o1144]='o0000;
mem_cp['o1145]='o0000;
mem_cp['o1146]='o0000;
mem_cp['o1147]='o0000;
mem_cp['o1150]='o0000;
mem_cp['o1151]='o0000;
mem_cp['o1152]='o0000;
mem_cp['o1153]='o0000;
mem_cp['o1154]='o0000;
mem_cp['o1155]='o0000;
mem_cp['o1156]='o0000;
mem_cp['o1157]='o0000;
mem_cp['o1160]='o0000;
mem_cp['o1161]='o0000;
mem_cp['o1162]='o0000;
mem_cp['o1163]='o0000;
mem_cp['o1164]='o0000;
mem_cp['o1165]='o0000;
mem_cp['o1166]='o0000;
mem_cp['o1167]='o0000;
mem_cp['o1170]='o0000;
mem_cp['o1171]='o0000;
mem_cp['o1172]='o0000;
mem_cp['o1173]='o0000;
mem_cp['o1174]='o0000;
mem_cp['o1175]='o0000;
mem_cp['o1176]='o0000;
mem_cp['o1177]='o0000;
mem_cp['o1200]='o0000;
mem_cp['o1201]='o0000;
mem_cp['o1202]='o0000;
mem_cp['o1203]='o0000;
mem_cp['o1204]='o0000;
mem_cp['o1205]='o0000;
mem_cp['o1206]='o0000;
mem_cp['o1207]='o0000;
mem_cp['o1210]='o0000;
mem_cp['o1211]='o0000;
mem_cp['o1212]='o0000;
mem_cp['o1213]='o0000;
mem_cp['o1214]='o0000;
mem_cp['o1215]='o0000;
mem_cp['o1216]='o0000;
mem_cp['o1217]='o0000;
mem_cp['o1220]='o0000;
mem_cp['o1221]='o0000;
mem_cp['o1222]='o0000;
mem_cp['o1223]='o0000;
mem_cp['o1224]='o0000;
mem_cp['o1225]='o0000;
mem_cp['o1226]='o0000;
mem_cp['o1227]='o0000;
mem_cp['o1230]='o0000;
mem_cp['o1231]='o0000;
mem_cp['o1232]='o0000;
mem_cp['o1233]='o0000;
mem_cp['o1234]='o0000;
mem_cp['o1235]='o0000;
mem_cp['o1236]='o0000;
mem_cp['o1237]='o0000;
mem_cp['o1240]='o0000;
mem_cp['o1241]='o0000;
mem_cp['o1242]='o0000;
mem_cp['o1243]='o0000;
mem_cp['o1244]='o0000;
mem_cp['o1245]='o0000;
mem_cp['o1246]='o0000;
mem_cp['o1247]='o0000;
mem_cp['o1250]='o0000;
mem_cp['o1251]='o0000;
mem_cp['o1252]='o0000;
mem_cp['o1253]='o0000;
mem_cp['o1254]='o0000;
mem_cp['o1255]='o0000;
mem_cp['o1256]='o0000;
mem_cp['o1257]='o0000;
mem_cp['o1260]='o0000;
mem_cp['o1261]='o0000;
mem_cp['o1262]='o0000;
mem_cp['o1263]='o0000;
mem_cp['o1264]='o0000;
mem_cp['o1265]='o0000;
mem_cp['o1266]='o0000;
mem_cp['o1267]='o0000;
mem_cp['o1270]='o0000;
mem_cp['o1271]='o0000;
mem_cp['o1272]='o0000;
mem_cp['o1273]='o0000;
mem_cp['o1274]='o0000;
mem_cp['o1275]='o0000;
mem_cp['o1276]='o0000;
mem_cp['o1277]='o0000;
mem_cp['o1300]='o0000;
mem_cp['o1301]='o0000;
mem_cp['o1302]='o0000;
mem_cp['o1303]='o0000;
mem_cp['o1304]='o0000;
mem_cp['o1305]='o0000;
mem_cp['o1306]='o0000;
mem_cp['o1307]='o0000;
mem_cp['o1310]='o0000;
mem_cp['o1311]='o0000;
mem_cp['o1312]='o0000;
mem_cp['o1313]='o0000;
mem_cp['o1314]='o0000;
mem_cp['o1315]='o0000;
mem_cp['o1316]='o0000;
mem_cp['o1317]='o0000;
mem_cp['o1320]='o0000;
mem_cp['o1321]='o0000;
mem_cp['o1322]='o0000;
mem_cp['o1323]='o0000;
mem_cp['o1324]='o0000;
mem_cp['o1325]='o0000;
mem_cp['o1326]='o0000;
mem_cp['o1327]='o0000;
mem_cp['o1330]='o0000;
mem_cp['o1331]='o0000;
mem_cp['o1332]='o0000;
mem_cp['o1333]='o0000;
mem_cp['o1334]='o0000;
mem_cp['o1335]='o0000;
mem_cp['o1336]='o0000;
mem_cp['o1337]='o0000;
mem_cp['o1340]='o0000;
mem_cp['o1341]='o0000;
mem_cp['o1342]='o0000;
mem_cp['o1343]='o0000;
mem_cp['o1344]='o0000;
mem_cp['o1345]='o0000;
mem_cp['o1346]='o0000;
mem_cp['o1347]='o0000;
mem_cp['o1350]='o0000;
mem_cp['o1351]='o0000;
mem_cp['o1352]='o0000;
mem_cp['o1353]='o0000;
mem_cp['o1354]='o0000;
mem_cp['o1355]='o0000;
mem_cp['o1356]='o0000;
mem_cp['o1357]='o0000;
mem_cp['o1360]='o0000;
mem_cp['o1361]='o0000;
mem_cp['o1362]='o0000;
mem_cp['o1363]='o0000;
mem_cp['o1364]='o0000;
mem_cp['o1365]='o0000;
mem_cp['o1366]='o0000;
mem_cp['o1367]='o0000;
mem_cp['o1370]='o0000;
mem_cp['o1371]='o0000;
mem_cp['o1372]='o0000;
mem_cp['o1373]='o0000;
mem_cp['o1374]='o0000;
mem_cp['o1375]='o0000;
mem_cp['o1376]='o0000;
mem_cp['o1377]='o0000;
mem_cp['o1400]='o0000;
mem_cp['o1401]='o0000;
mem_cp['o1402]='o0000;
mem_cp['o1403]='o0000;
mem_cp['o1404]='o0000;
mem_cp['o1405]='o0000;
mem_cp['o1406]='o0000;
mem_cp['o1407]='o0000;
mem_cp['o1410]='o0000;
mem_cp['o1411]='o0000;
mem_cp['o1412]='o0000;
mem_cp['o1413]='o0000;
mem_cp['o1414]='o0000;
mem_cp['o1415]='o0000;
mem_cp['o1416]='o0000;
mem_cp['o1417]='o0000;
mem_cp['o1420]='o0000;
mem_cp['o1421]='o0000;
mem_cp['o1422]='o0000;
mem_cp['o1423]='o0000;
mem_cp['o1424]='o0000;
mem_cp['o1425]='o0000;
mem_cp['o1426]='o0000;
mem_cp['o1427]='o0000;
mem_cp['o1430]='o0000;
mem_cp['o1431]='o0000;
mem_cp['o1432]='o0000;
mem_cp['o1433]='o0000;
mem_cp['o1434]='o0000;
mem_cp['o1435]='o0000;
mem_cp['o1436]='o0000;
mem_cp['o1437]='o0000;
mem_cp['o1440]='o0000;
mem_cp['o1441]='o0000;
mem_cp['o1442]='o0000;
mem_cp['o1443]='o0000;
mem_cp['o1444]='o0000;
mem_cp['o1445]='o0000;
mem_cp['o1446]='o0000;
mem_cp['o1447]='o0000;
mem_cp['o1450]='o0000;
mem_cp['o1451]='o0000;
mem_cp['o1452]='o0000;
mem_cp['o1453]='o0000;
mem_cp['o1454]='o0000;
mem_cp['o1455]='o0000;
mem_cp['o1456]='o0000;
mem_cp['o1457]='o0000;
mem_cp['o1460]='o0000;
mem_cp['o1461]='o0000;
mem_cp['o1462]='o0000;
mem_cp['o1463]='o0000;
mem_cp['o1464]='o0000;
mem_cp['o1465]='o0000;
mem_cp['o1466]='o0000;
mem_cp['o1467]='o0000;
mem_cp['o1470]='o0000;
mem_cp['o1471]='o0000;
mem_cp['o1472]='o0000;
mem_cp['o1473]='o0000;
mem_cp['o1474]='o0000;
mem_cp['o1475]='o0000;
mem_cp['o1476]='o0000;
mem_cp['o1477]='o0000;
mem_cp['o1500]='o0000;
mem_cp['o1501]='o0000;
mem_cp['o1502]='o0000;
mem_cp['o1503]='o0000;
mem_cp['o1504]='o0000;
mem_cp['o1505]='o0000;
mem_cp['o1506]='o0000;
mem_cp['o1507]='o0000;
mem_cp['o1510]='o0000;
mem_cp['o1511]='o0000;
mem_cp['o1512]='o0000;
mem_cp['o1513]='o0000;
mem_cp['o1514]='o0000;
mem_cp['o1515]='o0000;
mem_cp['o1516]='o0000;
mem_cp['o1517]='o0000;
mem_cp['o1520]='o0000;
mem_cp['o1521]='o0000;
mem_cp['o1522]='o0000;
mem_cp['o1523]='o0000;
mem_cp['o1524]='o0000;
mem_cp['o1525]='o0000;
mem_cp['o1526]='o0000;
mem_cp['o1527]='o0000;
mem_cp['o1530]='o0000;
mem_cp['o1531]='o0000;
mem_cp['o1532]='o0000;
mem_cp['o1533]='o0000;
mem_cp['o1534]='o0000;
mem_cp['o1535]='o0000;
mem_cp['o1536]='o0000;
mem_cp['o1537]='o0000;
mem_cp['o1540]='o0000;
mem_cp['o1541]='o0000;
mem_cp['o1542]='o0000;
mem_cp['o1543]='o0000;
mem_cp['o1544]='o0000;
mem_cp['o1545]='o0000;
mem_cp['o1546]='o0000;
mem_cp['o1547]='o0000;
mem_cp['o1550]='o0000;
mem_cp['o1551]='o0000;
mem_cp['o1552]='o0000;
mem_cp['o1553]='o0000;
mem_cp['o1554]='o0000;
mem_cp['o1555]='o0000;
mem_cp['o1556]='o0000;
mem_cp['o1557]='o0000;
mem_cp['o1560]='o0000;
mem_cp['o1561]='o0000;
mem_cp['o1562]='o0000;
mem_cp['o1563]='o0000;
mem_cp['o1564]='o0000;
mem_cp['o1565]='o0000;
mem_cp['o1566]='o0000;
mem_cp['o1567]='o0000;
mem_cp['o1570]='o0000;
mem_cp['o1571]='o0000;
mem_cp['o1572]='o0000;
mem_cp['o1573]='o0000;
mem_cp['o1574]='o0000;
mem_cp['o1575]='o0000;
mem_cp['o1576]='o0000;
mem_cp['o1577]='o0000;
mem_cp['o1600]='o0000;
mem_cp['o1601]='o0000;
mem_cp['o1602]='o0000;
mem_cp['o1603]='o0000;
mem_cp['o1604]='o0000;
mem_cp['o1605]='o0000;
mem_cp['o1606]='o0000;
mem_cp['o1607]='o0000;
mem_cp['o1610]='o0000;
mem_cp['o1611]='o0000;
mem_cp['o1612]='o0000;
mem_cp['o1613]='o0000;
mem_cp['o1614]='o0000;
mem_cp['o1615]='o0000;
mem_cp['o1616]='o0000;
mem_cp['o1617]='o0000;
mem_cp['o1620]='o0000;
mem_cp['o1621]='o0000;
mem_cp['o1622]='o0000;
mem_cp['o1623]='o0000;
mem_cp['o1624]='o0000;
mem_cp['o1625]='o0000;
mem_cp['o1626]='o0000;
mem_cp['o1627]='o0000;
mem_cp['o1630]='o0000;
mem_cp['o1631]='o0000;
mem_cp['o1632]='o0000;
mem_cp['o1633]='o0000;
mem_cp['o1634]='o0000;
mem_cp['o1635]='o0000;
mem_cp['o1636]='o0000;
mem_cp['o1637]='o0000;
mem_cp['o1640]='o0000;
mem_cp['o1641]='o0000;
mem_cp['o1642]='o0000;
mem_cp['o1643]='o0000;
mem_cp['o1644]='o0000;
mem_cp['o1645]='o0000;
mem_cp['o1646]='o0000;
mem_cp['o1647]='o0000;
mem_cp['o1650]='o0000;
mem_cp['o1651]='o0000;
mem_cp['o1652]='o0000;
mem_cp['o1653]='o0000;
mem_cp['o1654]='o0000;
mem_cp['o1655]='o0000;
mem_cp['o1656]='o0000;
mem_cp['o1657]='o0000;
mem_cp['o1660]='o0000;
mem_cp['o1661]='o0000;
mem_cp['o1662]='o0000;
mem_cp['o1663]='o0000;
mem_cp['o1664]='o0000;
mem_cp['o1665]='o0000;
mem_cp['o1666]='o0000;
mem_cp['o1667]='o0000;
mem_cp['o1670]='o0000;
mem_cp['o1671]='o0000;
mem_cp['o1672]='o0000;
mem_cp['o1673]='o0000;
mem_cp['o1674]='o0000;
mem_cp['o1675]='o0000;
mem_cp['o1676]='o0000;
mem_cp['o1677]='o0000;
mem_cp['o1700]='o0000;
mem_cp['o1701]='o0000;
mem_cp['o1702]='o0000;
mem_cp['o1703]='o0000;
mem_cp['o1704]='o0000;
mem_cp['o1705]='o0000;
mem_cp['o1706]='o0000;
mem_cp['o1707]='o0000;
mem_cp['o1710]='o0000;
mem_cp['o1711]='o0000;
mem_cp['o1712]='o0000;
mem_cp['o1713]='o0000;
mem_cp['o1714]='o0000;
mem_cp['o1715]='o0000;
mem_cp['o1716]='o0000;
mem_cp['o1717]='o0000;
mem_cp['o1720]='o0000;
mem_cp['o1721]='o0000;
mem_cp['o1722]='o0000;
mem_cp['o1723]='o0000;
mem_cp['o1724]='o0000;
mem_cp['o1725]='o0000;
mem_cp['o1726]='o0000;
mem_cp['o1727]='o0000;
mem_cp['o1730]='o0000;
mem_cp['o1731]='o0000;
mem_cp['o1732]='o0000;
mem_cp['o1733]='o0000;
mem_cp['o1734]='o0000;
mem_cp['o1735]='o0000;
mem_cp['o1736]='o0000;
mem_cp['o1737]='o0000;
mem_cp['o1740]='o0000;
mem_cp['o1741]='o0000;
mem_cp['o1742]='o0000;
mem_cp['o1743]='o0000;
mem_cp['o1744]='o0000;
mem_cp['o1745]='o0000;
mem_cp['o1746]='o0000;
mem_cp['o1747]='o0000;
mem_cp['o1750]='o0000;
mem_cp['o1751]='o0000;
mem_cp['o1752]='o0000;
mem_cp['o1753]='o0000;
mem_cp['o1754]='o0000;
mem_cp['o1755]='o0000;
mem_cp['o1756]='o0000;
mem_cp['o1757]='o0000;
mem_cp['o1760]='o0000;
mem_cp['o1761]='o0000;
mem_cp['o1762]='o0000;
mem_cp['o1763]='o0000;
mem_cp['o1764]='o0000;
mem_cp['o1765]='o0000;
mem_cp['o1766]='o0000;
mem_cp['o1767]='o0000;
mem_cp['o1770]='o0000;
mem_cp['o1771]='o0000;
mem_cp['o1772]='o0000;
mem_cp['o1773]='o0000;
mem_cp['o1774]='o0000;
mem_cp['o1775]='o0000;
mem_cp['o1776]='o0000;
mem_cp['o1777]='o0000;
mem_cp['o2000]='o0000;
mem_cp['o2001]='o0000;
mem_cp['o2002]='o0000;
mem_cp['o2003]='o0000;
mem_cp['o2004]='o0000;
mem_cp['o2005]='o0000;
mem_cp['o2006]='o0000;
mem_cp['o2007]='o0000;
mem_cp['o2010]='o0000;
mem_cp['o2011]='o0000;
mem_cp['o2012]='o0000;
mem_cp['o2013]='o0000;
mem_cp['o2014]='o0000;
mem_cp['o2015]='o0000;
mem_cp['o2016]='o0000;
mem_cp['o2017]='o0000;
mem_cp['o2020]='o0000;
mem_cp['o2021]='o0000;
mem_cp['o2022]='o0000;
mem_cp['o2023]='o0000;
mem_cp['o2024]='o0000;
mem_cp['o2025]='o0000;
mem_cp['o2026]='o0000;
mem_cp['o2027]='o0000;
mem_cp['o2030]='o0000;
mem_cp['o2031]='o0000;
mem_cp['o2032]='o0000;
mem_cp['o2033]='o0000;
mem_cp['o2034]='o0000;
mem_cp['o2035]='o0000;
mem_cp['o2036]='o0000;
mem_cp['o2037]='o0000;
mem_cp['o2040]='o0000;
mem_cp['o2041]='o0000;
mem_cp['o2042]='o0000;
mem_cp['o2043]='o0000;
mem_cp['o2044]='o0000;
mem_cp['o2045]='o0000;
mem_cp['o2046]='o0000;
mem_cp['o2047]='o0000;
mem_cp['o2050]='o0000;
mem_cp['o2051]='o0000;
mem_cp['o2052]='o0000;
mem_cp['o2053]='o0000;
mem_cp['o2054]='o0000;
mem_cp['o2055]='o0000;
mem_cp['o2056]='o0000;
mem_cp['o2057]='o0000;
mem_cp['o2060]='o0000;
mem_cp['o2061]='o0000;
mem_cp['o2062]='o0000;
mem_cp['o2063]='o0000;
mem_cp['o2064]='o0000;
mem_cp['o2065]='o0000;
mem_cp['o2066]='o0000;
mem_cp['o2067]='o0000;
mem_cp['o2070]='o0000;
mem_cp['o2071]='o0000;
mem_cp['o2072]='o0000;
mem_cp['o2073]='o0000;
mem_cp['o2074]='o0000;
mem_cp['o2075]='o0000;
mem_cp['o2076]='o0000;
mem_cp['o2077]='o0000;
mem_cp['o2100]='o0000;
mem_cp['o2101]='o0000;
mem_cp['o2102]='o0000;
mem_cp['o2103]='o0000;
mem_cp['o2104]='o0000;
mem_cp['o2105]='o0000;
mem_cp['o2106]='o0000;
mem_cp['o2107]='o0000;
mem_cp['o2110]='o0000;
mem_cp['o2111]='o0000;
mem_cp['o2112]='o0000;
mem_cp['o2113]='o0000;
mem_cp['o2114]='o0000;
mem_cp['o2115]='o0000;
mem_cp['o2116]='o0000;
mem_cp['o2117]='o0000;
mem_cp['o2120]='o0000;
mem_cp['o2121]='o0000;
mem_cp['o2122]='o0000;
mem_cp['o2123]='o0000;
mem_cp['o2124]='o0000;
mem_cp['o2125]='o0000;
mem_cp['o2126]='o0000;
mem_cp['o2127]='o0000;
mem_cp['o2130]='o0000;
mem_cp['o2131]='o0000;
mem_cp['o2132]='o0000;
mem_cp['o2133]='o0000;
mem_cp['o2134]='o0000;
mem_cp['o2135]='o0000;
mem_cp['o2136]='o0000;
mem_cp['o2137]='o0000;
mem_cp['o2140]='o0000;
mem_cp['o2141]='o0000;
mem_cp['o2142]='o0000;
mem_cp['o2143]='o0000;
mem_cp['o2144]='o0000;
mem_cp['o2145]='o0000;
mem_cp['o2146]='o0000;
mem_cp['o2147]='o0000;
mem_cp['o2150]='o0000;
mem_cp['o2151]='o0000;
mem_cp['o2152]='o0000;
mem_cp['o2153]='o0000;
mem_cp['o2154]='o0000;
mem_cp['o2155]='o0000;
mem_cp['o2156]='o0000;
mem_cp['o2157]='o0000;
mem_cp['o2160]='o0000;
mem_cp['o2161]='o0000;
mem_cp['o2162]='o0000;
mem_cp['o2163]='o0000;
mem_cp['o2164]='o0000;
mem_cp['o2165]='o0000;
mem_cp['o2166]='o0000;
mem_cp['o2167]='o0000;
mem_cp['o2170]='o0000;
mem_cp['o2171]='o0000;
mem_cp['o2172]='o0000;
mem_cp['o2173]='o0000;
mem_cp['o2174]='o0000;
mem_cp['o2175]='o0000;
mem_cp['o2176]='o0000;
mem_cp['o2177]='o0000;
mem_cp['o2200]='o0000;
mem_cp['o2201]='o0000;
mem_cp['o2202]='o0000;
mem_cp['o2203]='o0000;
mem_cp['o2204]='o0000;
mem_cp['o2205]='o0000;
mem_cp['o2206]='o0000;
mem_cp['o2207]='o0000;
mem_cp['o2210]='o0000;
mem_cp['o2211]='o0000;
mem_cp['o2212]='o0000;
mem_cp['o2213]='o0000;
mem_cp['o2214]='o0000;
mem_cp['o2215]='o0000;
mem_cp['o2216]='o0000;
mem_cp['o2217]='o0000;
mem_cp['o2220]='o0000;
mem_cp['o2221]='o0000;
mem_cp['o2222]='o0000;
mem_cp['o2223]='o0000;
mem_cp['o2224]='o0000;
mem_cp['o2225]='o0000;
mem_cp['o2226]='o0000;
mem_cp['o2227]='o0000;
mem_cp['o2230]='o0000;
mem_cp['o2231]='o0000;
mem_cp['o2232]='o0000;
mem_cp['o2233]='o0000;
mem_cp['o2234]='o0000;
mem_cp['o2235]='o0000;
mem_cp['o2236]='o0000;
mem_cp['o2237]='o0000;
mem_cp['o2240]='o0000;
mem_cp['o2241]='o0000;
mem_cp['o2242]='o0000;
mem_cp['o2243]='o0000;
mem_cp['o2244]='o0000;
mem_cp['o2245]='o0000;
mem_cp['o2246]='o0000;
mem_cp['o2247]='o0000;
mem_cp['o2250]='o0000;
mem_cp['o2251]='o0000;
mem_cp['o2252]='o0000;
mem_cp['o2253]='o0000;
mem_cp['o2254]='o0000;
mem_cp['o2255]='o0000;
mem_cp['o2256]='o0000;
mem_cp['o2257]='o0000;
mem_cp['o2260]='o0000;
mem_cp['o2261]='o0000;
mem_cp['o2262]='o0000;
mem_cp['o2263]='o0000;
mem_cp['o2264]='o0000;
mem_cp['o2265]='o0000;
mem_cp['o2266]='o0000;
mem_cp['o2267]='o0000;
mem_cp['o2270]='o0000;
mem_cp['o2271]='o0000;
mem_cp['o2272]='o0000;
mem_cp['o2273]='o0000;
mem_cp['o2274]='o0000;
mem_cp['o2275]='o0000;
mem_cp['o2276]='o0000;
mem_cp['o2277]='o0000;
mem_cp['o2300]='o0000;
mem_cp['o2301]='o0000;
mem_cp['o2302]='o0000;
mem_cp['o2303]='o0000;
mem_cp['o2304]='o0000;
mem_cp['o2305]='o0000;
mem_cp['o2306]='o0000;
mem_cp['o2307]='o0000;
mem_cp['o2310]='o0000;
mem_cp['o2311]='o0000;
mem_cp['o2312]='o0000;
mem_cp['o2313]='o0000;
mem_cp['o2314]='o0000;
mem_cp['o2315]='o0000;
mem_cp['o2316]='o0000;
mem_cp['o2317]='o0000;
mem_cp['o2320]='o0000;
mem_cp['o2321]='o0000;
mem_cp['o2322]='o0000;
mem_cp['o2323]='o0000;
mem_cp['o2324]='o0000;
mem_cp['o2325]='o0000;
mem_cp['o2326]='o0000;
mem_cp['o2327]='o0000;
mem_cp['o2330]='o0000;
mem_cp['o2331]='o0000;
mem_cp['o2332]='o0000;
mem_cp['o2333]='o0000;
mem_cp['o2334]='o0000;
mem_cp['o2335]='o0000;
mem_cp['o2336]='o0000;
mem_cp['o2337]='o0000;
mem_cp['o2340]='o0000;
mem_cp['o2341]='o0000;
mem_cp['o2342]='o0000;
mem_cp['o2343]='o0000;
mem_cp['o2344]='o0000;
mem_cp['o2345]='o0000;
mem_cp['o2346]='o0000;
mem_cp['o2347]='o0000;
mem_cp['o2350]='o0000;
mem_cp['o2351]='o0000;
mem_cp['o2352]='o0000;
mem_cp['o2353]='o0000;
mem_cp['o2354]='o0000;
mem_cp['o2355]='o0000;
mem_cp['o2356]='o0000;
mem_cp['o2357]='o0000;
mem_cp['o2360]='o0000;
mem_cp['o2361]='o0000;
mem_cp['o2362]='o0000;
mem_cp['o2363]='o0000;
mem_cp['o2364]='o0000;
mem_cp['o2365]='o0000;
mem_cp['o2366]='o0000;
mem_cp['o2367]='o0000;
mem_cp['o2370]='o0000;
mem_cp['o2371]='o0000;
mem_cp['o2372]='o0000;
mem_cp['o2373]='o0000;
mem_cp['o2374]='o0000;
mem_cp['o2375]='o0000;
mem_cp['o2376]='o0000;
mem_cp['o2377]='o0000;
mem_cp['o2400]='o0000;
mem_cp['o2401]='o0000;
mem_cp['o2402]='o0000;
mem_cp['o2403]='o0000;
mem_cp['o2404]='o0000;
mem_cp['o2405]='o0000;
mem_cp['o2406]='o0000;
mem_cp['o2407]='o0000;
mem_cp['o2410]='o0000;
mem_cp['o2411]='o0000;
mem_cp['o2412]='o0000;
mem_cp['o2413]='o0000;
mem_cp['o2414]='o0000;
mem_cp['o2415]='o0000;
mem_cp['o2416]='o0000;
mem_cp['o2417]='o0000;
mem_cp['o2420]='o0000;
mem_cp['o2421]='o0000;
mem_cp['o2422]='o0000;
mem_cp['o2423]='o0000;
mem_cp['o2424]='o0000;
mem_cp['o2425]='o0000;
mem_cp['o2426]='o0000;
mem_cp['o2427]='o0000;
mem_cp['o2430]='o0000;
mem_cp['o2431]='o0000;
mem_cp['o2432]='o0000;
mem_cp['o2433]='o0000;
mem_cp['o2434]='o0000;
mem_cp['o2435]='o0000;
mem_cp['o2436]='o0000;
mem_cp['o2437]='o0000;
mem_cp['o2440]='o0000;
mem_cp['o2441]='o0000;
mem_cp['o2442]='o0000;
mem_cp['o2443]='o0000;
mem_cp['o2444]='o0000;
mem_cp['o2445]='o0000;
mem_cp['o2446]='o0000;
mem_cp['o2447]='o0000;
mem_cp['o2450]='o0000;
mem_cp['o2451]='o0000;
mem_cp['o2452]='o0000;
mem_cp['o2453]='o0000;
mem_cp['o2454]='o0000;
mem_cp['o2455]='o0000;
mem_cp['o2456]='o0000;
mem_cp['o2457]='o0000;
mem_cp['o2460]='o0000;
mem_cp['o2461]='o0000;
mem_cp['o2462]='o0000;
mem_cp['o2463]='o0000;
mem_cp['o2464]='o0000;
mem_cp['o2465]='o0000;
mem_cp['o2466]='o0000;
mem_cp['o2467]='o0000;
mem_cp['o2470]='o0000;
mem_cp['o2471]='o0000;
mem_cp['o2472]='o0000;
mem_cp['o2473]='o0000;
mem_cp['o2474]='o0000;
mem_cp['o2475]='o0000;
mem_cp['o2476]='o0000;
mem_cp['o2477]='o0000;
mem_cp['o2500]='o0000;
mem_cp['o2501]='o0000;
mem_cp['o2502]='o0000;
mem_cp['o2503]='o0000;
mem_cp['o2504]='o0000;
mem_cp['o2505]='o0000;
mem_cp['o2506]='o0000;
mem_cp['o2507]='o0000;
mem_cp['o2510]='o0000;
mem_cp['o2511]='o0000;
mem_cp['o2512]='o0000;
mem_cp['o2513]='o0000;
mem_cp['o2514]='o0000;
mem_cp['o2515]='o0000;
mem_cp['o2516]='o0000;
mem_cp['o2517]='o0000;
mem_cp['o2520]='o0000;
mem_cp['o2521]='o0000;
mem_cp['o2522]='o0000;
mem_cp['o2523]='o0000;
mem_cp['o2524]='o0000;
mem_cp['o2525]='o0000;
mem_cp['o2526]='o0000;
mem_cp['o2527]='o0000;
mem_cp['o2530]='o0000;
mem_cp['o2531]='o0000;
mem_cp['o2532]='o0000;
mem_cp['o2533]='o0000;
mem_cp['o2534]='o0000;
mem_cp['o2535]='o0000;
mem_cp['o2536]='o0000;
mem_cp['o2537]='o0000;
mem_cp['o2540]='o0000;
mem_cp['o2541]='o0000;
mem_cp['o2542]='o0000;
mem_cp['o2543]='o0000;
mem_cp['o2544]='o0000;
mem_cp['o2545]='o0000;
mem_cp['o2546]='o0000;
mem_cp['o2547]='o0000;
mem_cp['o2550]='o0000;
mem_cp['o2551]='o0000;
mem_cp['o2552]='o0000;
mem_cp['o2553]='o0000;
mem_cp['o2554]='o0000;
mem_cp['o2555]='o0000;
mem_cp['o2556]='o0000;
mem_cp['o2557]='o0000;
mem_cp['o2560]='o0000;
mem_cp['o2561]='o0000;
mem_cp['o2562]='o0000;
mem_cp['o2563]='o0000;
mem_cp['o2564]='o0000;
mem_cp['o2565]='o0000;
mem_cp['o2566]='o0000;
mem_cp['o2567]='o0000;
mem_cp['o2570]='o0000;
mem_cp['o2571]='o0000;
mem_cp['o2572]='o0000;
mem_cp['o2573]='o0000;
mem_cp['o2574]='o0000;
mem_cp['o2575]='o0000;
mem_cp['o2576]='o0000;
mem_cp['o2577]='o0000;
mem_cp['o2600]='o0000;
mem_cp['o2601]='o0000;
mem_cp['o2602]='o0000;
mem_cp['o2603]='o0000;
mem_cp['o2604]='o0000;
mem_cp['o2605]='o0000;
mem_cp['o2606]='o0000;
mem_cp['o2607]='o0000;
mem_cp['o2610]='o0000;
mem_cp['o2611]='o0000;
mem_cp['o2612]='o0000;
mem_cp['o2613]='o0000;
mem_cp['o2614]='o0000;
mem_cp['o2615]='o0000;
mem_cp['o2616]='o0000;
mem_cp['o2617]='o0000;
mem_cp['o2620]='o0000;
mem_cp['o2621]='o0000;
mem_cp['o2622]='o0000;
mem_cp['o2623]='o0000;
mem_cp['o2624]='o0000;
mem_cp['o2625]='o0000;
mem_cp['o2626]='o0000;
mem_cp['o2627]='o0000;
mem_cp['o2630]='o0000;
mem_cp['o2631]='o0000;
mem_cp['o2632]='o0000;
mem_cp['o2633]='o0000;
mem_cp['o2634]='o0000;
mem_cp['o2635]='o0000;
mem_cp['o2636]='o0000;
mem_cp['o2637]='o0000;
mem_cp['o2640]='o0000;
mem_cp['o2641]='o0000;
mem_cp['o2642]='o0000;
mem_cp['o2643]='o0000;
mem_cp['o2644]='o0000;
mem_cp['o2645]='o0000;
mem_cp['o2646]='o0000;
mem_cp['o2647]='o0000;
mem_cp['o2650]='o0000;
mem_cp['o2651]='o0000;
mem_cp['o2652]='o0000;
mem_cp['o2653]='o0000;
mem_cp['o2654]='o0000;
mem_cp['o2655]='o0000;
mem_cp['o2656]='o0000;
mem_cp['o2657]='o0000;
mem_cp['o2660]='o0000;
mem_cp['o2661]='o0000;
mem_cp['o2662]='o0000;
mem_cp['o2663]='o0000;
mem_cp['o2664]='o0000;
mem_cp['o2665]='o0000;
mem_cp['o2666]='o0000;
mem_cp['o2667]='o0000;
mem_cp['o2670]='o0000;
mem_cp['o2671]='o0000;
mem_cp['o2672]='o0000;
mem_cp['o2673]='o0000;
mem_cp['o2674]='o0000;
mem_cp['o2675]='o0000;
mem_cp['o2676]='o0000;
mem_cp['o2677]='o0000;
mem_cp['o2700]='o0000;
mem_cp['o2701]='o0000;
mem_cp['o2702]='o0000;
mem_cp['o2703]='o0000;
mem_cp['o2704]='o0000;
mem_cp['o2705]='o0000;
mem_cp['o2706]='o0000;
mem_cp['o2707]='o0000;
mem_cp['o2710]='o0000;
mem_cp['o2711]='o0000;
mem_cp['o2712]='o0000;
mem_cp['o2713]='o0000;
mem_cp['o2714]='o0000;
mem_cp['o2715]='o0000;
mem_cp['o2716]='o0000;
mem_cp['o2717]='o0000;
mem_cp['o2720]='o0000;
mem_cp['o2721]='o0000;
mem_cp['o2722]='o0000;
mem_cp['o2723]='o0000;
mem_cp['o2724]='o0000;
mem_cp['o2725]='o0000;
mem_cp['o2726]='o0000;
mem_cp['o2727]='o0000;
mem_cp['o2730]='o0000;
mem_cp['o2731]='o0000;
mem_cp['o2732]='o0000;
mem_cp['o2733]='o0000;
mem_cp['o2734]='o0000;
mem_cp['o2735]='o0000;
mem_cp['o2736]='o0000;
mem_cp['o2737]='o0000;
mem_cp['o2740]='o0000;
mem_cp['o2741]='o0000;
mem_cp['o2742]='o0000;
mem_cp['o2743]='o0000;
mem_cp['o2744]='o0000;
mem_cp['o2745]='o0000;
mem_cp['o2746]='o0000;
mem_cp['o2747]='o0000;
mem_cp['o2750]='o0000;
mem_cp['o2751]='o0000;
mem_cp['o2752]='o0000;
mem_cp['o2753]='o0000;
mem_cp['o2754]='o0000;
mem_cp['o2755]='o0000;
mem_cp['o2756]='o0000;
mem_cp['o2757]='o0000;
mem_cp['o2760]='o0000;
mem_cp['o2761]='o0000;
mem_cp['o2762]='o0000;
mem_cp['o2763]='o0000;
mem_cp['o2764]='o0000;
mem_cp['o2765]='o0000;
mem_cp['o2766]='o0000;
mem_cp['o2767]='o0000;
mem_cp['o2770]='o0000;
mem_cp['o2771]='o0000;
mem_cp['o2772]='o0000;
mem_cp['o2773]='o0000;
mem_cp['o2774]='o0000;
mem_cp['o2775]='o0000;
mem_cp['o2776]='o0000;
mem_cp['o2777]='o0000;
mem_cp['o3000]='o0000;
mem_cp['o3001]='o0000;
mem_cp['o3002]='o0000;
mem_cp['o3003]='o0000;
mem_cp['o3004]='o0000;
mem_cp['o3005]='o0000;
mem_cp['o3006]='o0000;
mem_cp['o3007]='o0000;
mem_cp['o3010]='o0000;
mem_cp['o3011]='o0000;
mem_cp['o3012]='o0000;
mem_cp['o3013]='o0000;
mem_cp['o3014]='o0000;
mem_cp['o3015]='o0000;
mem_cp['o3016]='o0000;
mem_cp['o3017]='o0000;
mem_cp['o3020]='o0000;
mem_cp['o3021]='o0000;
mem_cp['o3022]='o0000;
mem_cp['o3023]='o0000;
mem_cp['o3024]='o0000;
mem_cp['o3025]='o0000;
mem_cp['o3026]='o0000;
mem_cp['o3027]='o0000;
mem_cp['o3030]='o0000;
mem_cp['o3031]='o0000;
mem_cp['o3032]='o0000;
mem_cp['o3033]='o0000;
mem_cp['o3034]='o0000;
mem_cp['o3035]='o0000;
mem_cp['o3036]='o0000;
mem_cp['o3037]='o0000;
mem_cp['o3040]='o0000;
mem_cp['o3041]='o0000;
mem_cp['o3042]='o0000;
mem_cp['o3043]='o0000;
mem_cp['o3044]='o0000;
mem_cp['o3045]='o0000;
mem_cp['o3046]='o0000;
mem_cp['o3047]='o0000;
mem_cp['o3050]='o0000;
mem_cp['o3051]='o0000;
mem_cp['o3052]='o0000;
mem_cp['o3053]='o0000;
mem_cp['o3054]='o0000;
mem_cp['o3055]='o0000;
mem_cp['o3056]='o0000;
mem_cp['o3057]='o0000;
mem_cp['o3060]='o0000;
mem_cp['o3061]='o0000;
mem_cp['o3062]='o0000;
mem_cp['o3063]='o0000;
mem_cp['o3064]='o0000;
mem_cp['o3065]='o0000;
mem_cp['o3066]='o0000;
mem_cp['o3067]='o0000;
mem_cp['o3070]='o0000;
mem_cp['o3071]='o0000;
mem_cp['o3072]='o0000;
mem_cp['o3073]='o0000;
mem_cp['o3074]='o0000;
mem_cp['o3075]='o0000;
mem_cp['o3076]='o0000;
mem_cp['o3077]='o0000;
mem_cp['o3100]='o0000;
mem_cp['o3101]='o0000;
mem_cp['o3102]='o0000;
mem_cp['o3103]='o0000;
mem_cp['o3104]='o0000;
mem_cp['o3105]='o0000;
mem_cp['o3106]='o0000;
mem_cp['o3107]='o0000;
mem_cp['o3110]='o0000;
mem_cp['o3111]='o0000;
mem_cp['o3112]='o0000;
mem_cp['o3113]='o0000;
mem_cp['o3114]='o0000;
mem_cp['o3115]='o0000;
mem_cp['o3116]='o0000;
mem_cp['o3117]='o0000;
mem_cp['o3120]='o0000;
mem_cp['o3121]='o0000;
mem_cp['o3122]='o0000;
mem_cp['o3123]='o0000;
mem_cp['o3124]='o0000;
mem_cp['o3125]='o0000;
mem_cp['o3126]='o0000;
mem_cp['o3127]='o0000;
mem_cp['o3130]='o0000;
mem_cp['o3131]='o0000;
mem_cp['o3132]='o0000;
mem_cp['o3133]='o0000;
mem_cp['o3134]='o0000;
mem_cp['o3135]='o0000;
mem_cp['o3136]='o0000;
mem_cp['o3137]='o0000;
mem_cp['o3140]='o0000;
mem_cp['o3141]='o0000;
mem_cp['o3142]='o0000;
mem_cp['o3143]='o0000;
mem_cp['o3144]='o0000;
mem_cp['o3145]='o0000;
mem_cp['o3146]='o0000;
mem_cp['o3147]='o0000;
mem_cp['o3150]='o0000;
mem_cp['o3151]='o0000;
mem_cp['o3152]='o0000;
mem_cp['o3153]='o0000;
mem_cp['o3154]='o0000;
mem_cp['o3155]='o0000;
mem_cp['o3156]='o0000;
mem_cp['o3157]='o0000;
mem_cp['o3160]='o0000;
mem_cp['o3161]='o0000;
mem_cp['o3162]='o0000;
mem_cp['o3163]='o0000;
mem_cp['o3164]='o0000;
mem_cp['o3165]='o0000;
mem_cp['o3166]='o0000;
mem_cp['o3167]='o0000;
mem_cp['o3170]='o0000;
mem_cp['o3171]='o0000;
mem_cp['o3172]='o0000;
mem_cp['o3173]='o0000;
mem_cp['o3174]='o0000;
mem_cp['o3175]='o0000;
mem_cp['o3176]='o0000;
mem_cp['o3177]='o0000;
mem_cp['o3200]='o0000;
mem_cp['o3201]='o0000;
mem_cp['o3202]='o0000;
mem_cp['o3203]='o0000;
mem_cp['o3204]='o0000;
mem_cp['o3205]='o0000;
mem_cp['o3206]='o0000;
mem_cp['o3207]='o0000;
mem_cp['o3210]='o0000;
mem_cp['o3211]='o0000;
mem_cp['o3212]='o0000;
mem_cp['o3213]='o0000;
mem_cp['o3214]='o0000;
mem_cp['o3215]='o0000;
mem_cp['o3216]='o0000;
mem_cp['o3217]='o0000;
mem_cp['o3220]='o0000;
mem_cp['o3221]='o0000;
mem_cp['o3222]='o0000;
mem_cp['o3223]='o0000;
mem_cp['o3224]='o0000;
mem_cp['o3225]='o0000;
mem_cp['o3226]='o0000;
mem_cp['o3227]='o0000;
mem_cp['o3230]='o0000;
mem_cp['o3231]='o0000;
mem_cp['o3232]='o0000;
mem_cp['o3233]='o0000;
mem_cp['o3234]='o0000;
mem_cp['o3235]='o0000;
mem_cp['o3236]='o0000;
mem_cp['o3237]='o0000;
mem_cp['o3240]='o0000;
mem_cp['o3241]='o0000;
mem_cp['o3242]='o0000;
mem_cp['o3243]='o0000;
mem_cp['o3244]='o0000;
mem_cp['o3245]='o0000;
mem_cp['o3246]='o0000;
mem_cp['o3247]='o0000;
mem_cp['o3250]='o0000;
mem_cp['o3251]='o0000;
mem_cp['o3252]='o0000;
mem_cp['o3253]='o0000;
mem_cp['o3254]='o0000;
mem_cp['o3255]='o0000;
mem_cp['o3256]='o0000;
mem_cp['o3257]='o0000;
mem_cp['o3260]='o0000;
mem_cp['o3261]='o0000;
mem_cp['o3262]='o0000;
mem_cp['o3263]='o0000;
mem_cp['o3264]='o0000;
mem_cp['o3265]='o0000;
mem_cp['o3266]='o0000;
mem_cp['o3267]='o0000;
mem_cp['o3270]='o0000;
mem_cp['o3271]='o0000;
mem_cp['o3272]='o0000;
mem_cp['o3273]='o0000;
mem_cp['o3274]='o0000;
mem_cp['o3275]='o0000;
mem_cp['o3276]='o0000;
mem_cp['o3277]='o0000;
mem_cp['o3300]='o0000;
mem_cp['o3301]='o0000;
mem_cp['o3302]='o0000;
mem_cp['o3303]='o0000;
mem_cp['o3304]='o0000;
mem_cp['o3305]='o0000;
mem_cp['o3306]='o0000;
mem_cp['o3307]='o0000;
mem_cp['o3310]='o0000;
mem_cp['o3311]='o0000;
mem_cp['o3312]='o0000;
mem_cp['o3313]='o0000;
mem_cp['o3314]='o0000;
mem_cp['o3315]='o0000;
mem_cp['o3316]='o0000;
mem_cp['o3317]='o0000;
mem_cp['o3320]='o0000;
mem_cp['o3321]='o0000;
mem_cp['o3322]='o0000;
mem_cp['o3323]='o0000;
mem_cp['o3324]='o0000;
mem_cp['o3325]='o0000;
mem_cp['o3326]='o0000;
mem_cp['o3327]='o0000;
mem_cp['o3330]='o0000;
mem_cp['o3331]='o0000;
mem_cp['o3332]='o0000;
mem_cp['o3333]='o0000;
mem_cp['o3334]='o0000;
mem_cp['o3335]='o0000;
mem_cp['o3336]='o0000;
mem_cp['o3337]='o0000;
mem_cp['o3340]='o0000;
mem_cp['o3341]='o0000;
mem_cp['o3342]='o0000;
mem_cp['o3343]='o0000;
mem_cp['o3344]='o0000;
mem_cp['o3345]='o0000;
mem_cp['o3346]='o0000;
mem_cp['o3347]='o0000;
mem_cp['o3350]='o0000;
mem_cp['o3351]='o0000;
mem_cp['o3352]='o0000;
mem_cp['o3353]='o0000;
mem_cp['o3354]='o0000;
mem_cp['o3355]='o0000;
mem_cp['o3356]='o0000;
mem_cp['o3357]='o0000;
mem_cp['o3360]='o0000;
mem_cp['o3361]='o0000;
mem_cp['o3362]='o0000;
mem_cp['o3363]='o0000;
mem_cp['o3364]='o0000;
mem_cp['o3365]='o0000;
mem_cp['o3366]='o0000;
mem_cp['o3367]='o0000;
mem_cp['o3370]='o0000;
mem_cp['o3371]='o0000;
mem_cp['o3372]='o0000;
mem_cp['o3373]='o0000;
mem_cp['o3374]='o0000;
mem_cp['o3375]='o0000;
mem_cp['o3376]='o0000;
mem_cp['o3377]='o0000;
mem_cp['o3400]='o0000;
mem_cp['o3401]='o0000;
mem_cp['o3402]='o0000;
mem_cp['o3403]='o0000;
mem_cp['o3404]='o0000;
mem_cp['o3405]='o0000;
mem_cp['o3406]='o0000;
mem_cp['o3407]='o0000;
mem_cp['o3410]='o0000;
mem_cp['o3411]='o0000;
mem_cp['o3412]='o0000;
mem_cp['o3413]='o0000;
mem_cp['o3414]='o0000;
mem_cp['o3415]='o0000;
mem_cp['o3416]='o0000;
mem_cp['o3417]='o0000;
mem_cp['o3420]='o0000;
mem_cp['o3421]='o0000;
mem_cp['o3422]='o0000;
mem_cp['o3423]='o0000;
mem_cp['o3424]='o0000;
mem_cp['o3425]='o0000;
mem_cp['o3426]='o0000;
mem_cp['o3427]='o0000;
mem_cp['o3430]='o0000;
mem_cp['o3431]='o0000;
mem_cp['o3432]='o0000;
mem_cp['o3433]='o0000;
mem_cp['o3434]='o0000;
mem_cp['o3435]='o0000;
mem_cp['o3436]='o0000;
mem_cp['o3437]='o0000;
mem_cp['o3440]='o0000;
mem_cp['o3441]='o0000;
mem_cp['o3442]='o0000;
mem_cp['o3443]='o0000;
mem_cp['o3444]='o0000;
mem_cp['o3445]='o0000;
mem_cp['o3446]='o0000;
mem_cp['o3447]='o0000;
mem_cp['o3450]='o0000;
mem_cp['o3451]='o0000;
mem_cp['o3452]='o0000;
mem_cp['o3453]='o0000;
mem_cp['o3454]='o0000;
mem_cp['o3455]='o0000;
mem_cp['o3456]='o0000;
mem_cp['o3457]='o0000;
mem_cp['o3460]='o0000;
mem_cp['o3461]='o0000;
mem_cp['o3462]='o0000;
mem_cp['o3463]='o0000;
mem_cp['o3464]='o0000;
mem_cp['o3465]='o0000;
mem_cp['o3466]='o0000;
mem_cp['o3467]='o0000;
mem_cp['o3470]='o0000;
mem_cp['o3471]='o0000;
mem_cp['o3472]='o0000;
mem_cp['o3473]='o0000;
mem_cp['o3474]='o0000;
mem_cp['o3475]='o0000;
mem_cp['o3476]='o0000;
mem_cp['o3477]='o0000;
mem_cp['o3500]='o0000;
mem_cp['o3501]='o0000;
mem_cp['o3502]='o0000;
mem_cp['o3503]='o0000;
mem_cp['o3504]='o0000;
mem_cp['o3505]='o0000;
mem_cp['o3506]='o0000;
mem_cp['o3507]='o0000;
mem_cp['o3510]='o0000;
mem_cp['o3511]='o0000;
mem_cp['o3512]='o0000;
mem_cp['o3513]='o0000;
mem_cp['o3514]='o0000;
mem_cp['o3515]='o0000;
mem_cp['o3516]='o0000;
mem_cp['o3517]='o0000;
mem_cp['o3520]='o0000;
mem_cp['o3521]='o0000;
mem_cp['o3522]='o0000;
mem_cp['o3523]='o0000;
mem_cp['o3524]='o0000;
mem_cp['o3525]='o0000;
mem_cp['o3526]='o0000;
mem_cp['o3527]='o0000;
mem_cp['o3530]='o0000;
mem_cp['o3531]='o0000;
mem_cp['o3532]='o0000;
mem_cp['o3533]='o0000;
mem_cp['o3534]='o0000;
mem_cp['o3535]='o0000;
mem_cp['o3536]='o0000;
mem_cp['o3537]='o0000;
mem_cp['o3540]='o0000;
mem_cp['o3541]='o0000;
mem_cp['o3542]='o0000;
mem_cp['o3543]='o0000;
mem_cp['o3544]='o0000;
mem_cp['o3545]='o0000;
mem_cp['o3546]='o0000;
mem_cp['o3547]='o0000;
mem_cp['o3550]='o0000;
mem_cp['o3551]='o0000;
mem_cp['o3552]='o0000;
mem_cp['o3553]='o0000;
mem_cp['o3554]='o0000;
mem_cp['o3555]='o0000;
mem_cp['o3556]='o0000;
mem_cp['o3557]='o0000;
mem_cp['o3560]='o0000;
mem_cp['o3561]='o0000;
mem_cp['o3562]='o0000;
mem_cp['o3563]='o0000;
mem_cp['o3564]='o0000;
mem_cp['o3565]='o0000;
mem_cp['o3566]='o0000;
mem_cp['o3567]='o0000;
mem_cp['o3570]='o0000;
mem_cp['o3571]='o0000;
mem_cp['o3572]='o0000;
mem_cp['o3573]='o0000;
mem_cp['o3574]='o0000;
mem_cp['o3575]='o0000;
mem_cp['o3576]='o0000;
mem_cp['o3577]='o0000;
mem_cp['o3600]='o0000;
mem_cp['o3601]='o0000;
mem_cp['o3602]='o0000;
mem_cp['o3603]='o0000;
mem_cp['o3604]='o0000;
mem_cp['o3605]='o0000;
mem_cp['o3606]='o0000;
mem_cp['o3607]='o0000;
mem_cp['o3610]='o0000;
mem_cp['o3611]='o0000;
mem_cp['o3612]='o0000;
mem_cp['o3613]='o0000;
mem_cp['o3614]='o0000;
mem_cp['o3615]='o0000;
mem_cp['o3616]='o0000;
mem_cp['o3617]='o0000;
mem_cp['o3620]='o0000;
mem_cp['o3621]='o0000;
mem_cp['o3622]='o0000;
mem_cp['o3623]='o0000;
mem_cp['o3624]='o0000;
mem_cp['o3625]='o0000;
mem_cp['o3626]='o0000;
mem_cp['o3627]='o0000;
mem_cp['o3630]='o0000;
mem_cp['o3631]='o0000;
mem_cp['o3632]='o0000;
mem_cp['o3633]='o0000;
mem_cp['o3634]='o0000;
mem_cp['o3635]='o0000;
mem_cp['o3636]='o0000;
mem_cp['o3637]='o0000;
mem_cp['o3640]='o0000;
mem_cp['o3641]='o0000;
mem_cp['o3642]='o0000;
mem_cp['o3643]='o0000;
mem_cp['o3644]='o0000;
mem_cp['o3645]='o0000;
mem_cp['o3646]='o0000;
mem_cp['o3647]='o0000;
mem_cp['o3650]='o0000;
mem_cp['o3651]='o0000;
mem_cp['o3652]='o0000;
mem_cp['o3653]='o0000;
mem_cp['o3654]='o0000;
mem_cp['o3655]='o0000;
mem_cp['o3656]='o0000;
mem_cp['o3657]='o0000;
mem_cp['o3660]='o0000;
mem_cp['o3661]='o0000;
mem_cp['o3662]='o0000;
mem_cp['o3663]='o0000;
mem_cp['o3664]='o0000;
mem_cp['o3665]='o0000;
mem_cp['o3666]='o0000;
mem_cp['o3667]='o0000;
mem_cp['o3670]='o0000;
mem_cp['o3671]='o0000;
mem_cp['o3672]='o0000;
mem_cp['o3673]='o0000;
mem_cp['o3674]='o0000;
mem_cp['o3675]='o0000;
mem_cp['o3676]='o0000;
mem_cp['o3677]='o0000;
mem_cp['o3700]='o0000;
mem_cp['o3701]='o0000;
mem_cp['o3702]='o0000;
mem_cp['o3703]='o0000;
mem_cp['o3704]='o0000;
mem_cp['o3705]='o0000;
mem_cp['o3706]='o0000;
mem_cp['o3707]='o0000;
mem_cp['o3710]='o0000;
mem_cp['o3711]='o0000;
mem_cp['o3712]='o0000;
mem_cp['o3713]='o0000;
mem_cp['o3714]='o0000;
mem_cp['o3715]='o0000;
mem_cp['o3716]='o0000;
mem_cp['o3717]='o0000;
mem_cp['o3720]='o0000;
mem_cp['o3721]='o0000;
mem_cp['o3722]='o0000;
mem_cp['o3723]='o0000;
mem_cp['o3724]='o0000;
mem_cp['o3725]='o0000;
mem_cp['o3726]='o0000;
mem_cp['o3727]='o0000;
mem_cp['o3730]='o0000;
mem_cp['o3731]='o0000;
mem_cp['o3732]='o0000;
mem_cp['o3733]='o0000;
mem_cp['o3734]='o0000;
mem_cp['o3735]='o0000;
mem_cp['o3736]='o0000;
mem_cp['o3737]='o0000;
mem_cp['o3740]='o0000;
mem_cp['o3741]='o0000;
mem_cp['o3742]='o0000;
mem_cp['o3743]='o0000;
mem_cp['o3744]='o0000;
mem_cp['o3745]='o0000;
mem_cp['o3746]='o0000;
mem_cp['o3747]='o0000;
mem_cp['o3750]='o0000;
mem_cp['o3751]='o0000;
mem_cp['o3752]='o0000;
mem_cp['o3753]='o0000;
mem_cp['o3754]='o0000;
mem_cp['o3755]='o0000;
mem_cp['o3756]='o0000;
mem_cp['o3757]='o0000;
mem_cp['o3760]='o0000;
mem_cp['o3761]='o0000;
mem_cp['o3762]='o0000;
mem_cp['o3763]='o0000;
mem_cp['o3764]='o0000;
mem_cp['o3765]='o0000;
mem_cp['o3766]='o0000;
mem_cp['o3767]='o0000;
mem_cp['o3770]='o0000;
mem_cp['o3771]='o0000;
mem_cp['o3772]='o0000;
mem_cp['o3773]='o0000;
mem_cp['o3774]='o0000;
mem_cp['o3775]='o0000;
mem_cp['o3776]='o0000;
mem_cp['o3777]='o0000;
mem_cp['o4000]='o0000;
mem_cp['o4001]='o0000;
mem_cp['o4002]='o0000;
mem_cp['o4003]='o0000;
mem_cp['o4004]='o0000;
mem_cp['o4005]='o0000;
mem_cp['o4006]='o0000;
mem_cp['o4007]='o0000;
mem_cp['o4010]='o0000;
mem_cp['o4011]='o0000;
mem_cp['o4012]='o0000;
mem_cp['o4013]='o0000;
mem_cp['o4014]='o0000;
mem_cp['o4015]='o0000;
mem_cp['o4016]='o0000;
mem_cp['o4017]='o0000;
mem_cp['o4020]='o0000;
mem_cp['o4021]='o0000;
mem_cp['o4022]='o0000;
mem_cp['o4023]='o0000;
mem_cp['o4024]='o0000;
mem_cp['o4025]='o0000;
mem_cp['o4026]='o0000;
mem_cp['o4027]='o0000;
mem_cp['o4030]='o0000;
mem_cp['o4031]='o0000;
mem_cp['o4032]='o0000;
mem_cp['o4033]='o0000;
mem_cp['o4034]='o0000;
mem_cp['o4035]='o0000;
mem_cp['o4036]='o0000;
mem_cp['o4037]='o0000;
mem_cp['o4040]='o0000;
mem_cp['o4041]='o0000;
mem_cp['o4042]='o0000;
mem_cp['o4043]='o0000;
mem_cp['o4044]='o0000;
mem_cp['o4045]='o0000;
mem_cp['o4046]='o0000;
mem_cp['o4047]='o0000;
mem_cp['o4050]='o0000;
mem_cp['o4051]='o0000;
mem_cp['o4052]='o0000;
mem_cp['o4053]='o0000;
mem_cp['o4054]='o0000;
mem_cp['o4055]='o0000;
mem_cp['o4056]='o0000;
mem_cp['o4057]='o0000;
mem_cp['o4060]='o0000;
mem_cp['o4061]='o0000;
mem_cp['o4062]='o0000;
mem_cp['o4063]='o0000;
mem_cp['o4064]='o0000;
mem_cp['o4065]='o0000;
mem_cp['o4066]='o0000;
mem_cp['o4067]='o0000;
mem_cp['o4070]='o0000;
mem_cp['o4071]='o0000;
mem_cp['o4072]='o0000;
mem_cp['o4073]='o0000;
mem_cp['o4074]='o0000;
mem_cp['o4075]='o0000;
mem_cp['o4076]='o0000;
mem_cp['o4077]='o0000;
mem_cp['o4100]='o0000;
mem_cp['o4101]='o0000;
mem_cp['o4102]='o0000;
mem_cp['o4103]='o0000;
mem_cp['o4104]='o0000;
mem_cp['o4105]='o0000;
mem_cp['o4106]='o0000;
mem_cp['o4107]='o0000;
mem_cp['o4110]='o0000;
mem_cp['o4111]='o0000;
mem_cp['o4112]='o0000;
mem_cp['o4113]='o0000;
mem_cp['o4114]='o0000;
mem_cp['o4115]='o0000;
mem_cp['o4116]='o0000;
mem_cp['o4117]='o0000;
mem_cp['o4120]='o0000;
mem_cp['o4121]='o0000;
mem_cp['o4122]='o0000;
mem_cp['o4123]='o0000;
mem_cp['o4124]='o0000;
mem_cp['o4125]='o0000;
mem_cp['o4126]='o0000;
mem_cp['o4127]='o0000;
mem_cp['o4130]='o0000;
mem_cp['o4131]='o0000;
mem_cp['o4132]='o0000;
mem_cp['o4133]='o0000;
mem_cp['o4134]='o0000;
mem_cp['o4135]='o0000;
mem_cp['o4136]='o0000;
mem_cp['o4137]='o0000;
mem_cp['o4140]='o0000;
mem_cp['o4141]='o0000;
mem_cp['o4142]='o0000;
mem_cp['o4143]='o0000;
mem_cp['o4144]='o0000;
mem_cp['o4145]='o0000;
mem_cp['o4146]='o0000;
mem_cp['o4147]='o0000;
mem_cp['o4150]='o0000;
mem_cp['o4151]='o0000;
mem_cp['o4152]='o0000;
mem_cp['o4153]='o0000;
mem_cp['o4154]='o0000;
mem_cp['o4155]='o0000;
mem_cp['o4156]='o0000;
mem_cp['o4157]='o0000;
mem_cp['o4160]='o0000;
mem_cp['o4161]='o0000;
mem_cp['o4162]='o0000;
mem_cp['o4163]='o0000;
mem_cp['o4164]='o0000;
mem_cp['o4165]='o0000;
mem_cp['o4166]='o0000;
mem_cp['o4167]='o0000;
mem_cp['o4170]='o0000;
mem_cp['o4171]='o0000;
mem_cp['o4172]='o0000;
mem_cp['o4173]='o0000;
mem_cp['o4174]='o0000;
mem_cp['o4175]='o0000;
mem_cp['o4176]='o0000;
mem_cp['o4177]='o0000;
mem_cp['o4200]='o0000;
mem_cp['o4201]='o0000;
mem_cp['o4202]='o0000;
mem_cp['o4203]='o0000;
mem_cp['o4204]='o0000;
mem_cp['o4205]='o0000;
mem_cp['o4206]='o0000;
mem_cp['o4207]='o0000;
mem_cp['o4210]='o0000;
mem_cp['o4211]='o0000;
mem_cp['o4212]='o0000;
mem_cp['o4213]='o0000;
mem_cp['o4214]='o0000;
mem_cp['o4215]='o0000;
mem_cp['o4216]='o0000;
mem_cp['o4217]='o0000;
mem_cp['o4220]='o0000;
mem_cp['o4221]='o0000;
mem_cp['o4222]='o0000;
mem_cp['o4223]='o0000;
mem_cp['o4224]='o0000;
mem_cp['o4225]='o0000;
mem_cp['o4226]='o0000;
mem_cp['o4227]='o0000;
mem_cp['o4230]='o0000;
mem_cp['o4231]='o0000;
mem_cp['o4232]='o0000;
mem_cp['o4233]='o0000;
mem_cp['o4234]='o0000;
mem_cp['o4235]='o0000;
mem_cp['o4236]='o0000;
mem_cp['o4237]='o0000;
mem_cp['o4240]='o0000;
mem_cp['o4241]='o0000;
mem_cp['o4242]='o0000;
mem_cp['o4243]='o0000;
mem_cp['o4244]='o0000;
mem_cp['o4245]='o0000;
mem_cp['o4246]='o0000;
mem_cp['o4247]='o0000;
mem_cp['o4250]='o0000;
mem_cp['o4251]='o0000;
mem_cp['o4252]='o0000;
mem_cp['o4253]='o0000;
mem_cp['o4254]='o0000;
mem_cp['o4255]='o0000;
mem_cp['o4256]='o0000;
mem_cp['o4257]='o0000;
mem_cp['o4260]='o0000;
mem_cp['o4261]='o0000;
mem_cp['o4262]='o0000;
mem_cp['o4263]='o0000;
mem_cp['o4264]='o0000;
mem_cp['o4265]='o0000;
mem_cp['o4266]='o0000;
mem_cp['o4267]='o0000;
mem_cp['o4270]='o0000;
mem_cp['o4271]='o0000;
mem_cp['o4272]='o0000;
mem_cp['o4273]='o0000;
mem_cp['o4274]='o0000;
mem_cp['o4275]='o0000;
mem_cp['o4276]='o0000;
mem_cp['o4277]='o0000;
mem_cp['o4300]='o0000;
mem_cp['o4301]='o0000;
mem_cp['o4302]='o0000;
mem_cp['o4303]='o0000;
mem_cp['o4304]='o0000;
mem_cp['o4305]='o0000;
mem_cp['o4306]='o0000;
mem_cp['o4307]='o0000;
mem_cp['o4310]='o0000;
mem_cp['o4311]='o0000;
mem_cp['o4312]='o0000;
mem_cp['o4313]='o0000;
mem_cp['o4314]='o0000;
mem_cp['o4315]='o0000;
mem_cp['o4316]='o0000;
mem_cp['o4317]='o0000;
mem_cp['o4320]='o0000;
mem_cp['o4321]='o0000;
mem_cp['o4322]='o0000;
mem_cp['o4323]='o0000;
mem_cp['o4324]='o0000;
mem_cp['o4325]='o0000;
mem_cp['o4326]='o0000;
mem_cp['o4327]='o0000;
mem_cp['o4330]='o0000;
mem_cp['o4331]='o0000;
mem_cp['o4332]='o0000;
mem_cp['o4333]='o0000;
mem_cp['o4334]='o0000;
mem_cp['o4335]='o0000;
mem_cp['o4336]='o0000;
mem_cp['o4337]='o0000;
mem_cp['o4340]='o0000;
mem_cp['o4341]='o0000;
mem_cp['o4342]='o0000;
mem_cp['o4343]='o0000;
mem_cp['o4344]='o0000;
mem_cp['o4345]='o0000;
mem_cp['o4346]='o0000;
mem_cp['o4347]='o0000;
mem_cp['o4350]='o0000;
mem_cp['o4351]='o0000;
mem_cp['o4352]='o0000;
mem_cp['o4353]='o0000;
mem_cp['o4354]='o0000;
mem_cp['o4355]='o0000;
mem_cp['o4356]='o0000;
mem_cp['o4357]='o0000;
mem_cp['o4360]='o0000;
mem_cp['o4361]='o0000;
mem_cp['o4362]='o0000;
mem_cp['o4363]='o0000;
mem_cp['o4364]='o0000;
mem_cp['o4365]='o0000;
mem_cp['o4366]='o0000;
mem_cp['o4367]='o0000;
mem_cp['o4370]='o0000;
mem_cp['o4371]='o0000;
mem_cp['o4372]='o0000;
mem_cp['o4373]='o0000;
mem_cp['o4374]='o0000;
mem_cp['o4375]='o0000;
mem_cp['o4376]='o0000;
mem_cp['o4377]='o0000;
mem_cp['o4400]='o0000;
mem_cp['o4401]='o0000;
mem_cp['o4402]='o0000;
mem_cp['o4403]='o0000;
mem_cp['o4404]='o0000;
mem_cp['o4405]='o0000;
mem_cp['o4406]='o0000;
mem_cp['o4407]='o0000;
mem_cp['o4410]='o0000;
mem_cp['o4411]='o0000;
mem_cp['o4412]='o0000;
mem_cp['o4413]='o0000;
mem_cp['o4414]='o0000;
mem_cp['o4415]='o0000;
mem_cp['o4416]='o0000;
mem_cp['o4417]='o0000;
mem_cp['o4420]='o0000;
mem_cp['o4421]='o0000;
mem_cp['o4422]='o0000;
mem_cp['o4423]='o0000;
mem_cp['o4424]='o0000;
mem_cp['o4425]='o0000;
mem_cp['o4426]='o0000;
mem_cp['o4427]='o0000;
mem_cp['o4430]='o0000;
mem_cp['o4431]='o0000;
mem_cp['o4432]='o0000;
mem_cp['o4433]='o0000;
mem_cp['o4434]='o0000;
mem_cp['o4435]='o0000;
mem_cp['o4436]='o0000;
mem_cp['o4437]='o0000;
mem_cp['o4440]='o0000;
mem_cp['o4441]='o0000;
mem_cp['o4442]='o0000;
mem_cp['o4443]='o0000;
mem_cp['o4444]='o0000;
mem_cp['o4445]='o0000;
mem_cp['o4446]='o0000;
mem_cp['o4447]='o0000;
mem_cp['o4450]='o0000;
mem_cp['o4451]='o0000;
mem_cp['o4452]='o0000;
mem_cp['o4453]='o0000;
mem_cp['o4454]='o0000;
mem_cp['o4455]='o0000;
mem_cp['o4456]='o0000;
mem_cp['o4457]='o0000;
mem_cp['o4460]='o0000;
mem_cp['o4461]='o0000;
mem_cp['o4462]='o0000;
mem_cp['o4463]='o0000;
mem_cp['o4464]='o0000;
mem_cp['o4465]='o0000;
mem_cp['o4466]='o0000;
mem_cp['o4467]='o0000;
mem_cp['o4470]='o0000;
mem_cp['o4471]='o0000;
mem_cp['o4472]='o0000;
mem_cp['o4473]='o0000;
mem_cp['o4474]='o0000;
mem_cp['o4475]='o0000;
mem_cp['o4476]='o0000;
mem_cp['o4477]='o0000;
mem_cp['o4500]='o0000;
mem_cp['o4501]='o0000;
mem_cp['o4502]='o0000;
mem_cp['o4503]='o0000;
mem_cp['o4504]='o0000;
mem_cp['o4505]='o0000;
mem_cp['o4506]='o0000;
mem_cp['o4507]='o0000;
mem_cp['o4510]='o0000;
mem_cp['o4511]='o0000;
mem_cp['o4512]='o0000;
mem_cp['o4513]='o0000;
mem_cp['o4514]='o0000;
mem_cp['o4515]='o0000;
mem_cp['o4516]='o0000;
mem_cp['o4517]='o0000;
mem_cp['o4520]='o0000;
mem_cp['o4521]='o0000;
mem_cp['o4522]='o0000;
mem_cp['o4523]='o0000;
mem_cp['o4524]='o0000;
mem_cp['o4525]='o0000;
mem_cp['o4526]='o0000;
mem_cp['o4527]='o0000;
mem_cp['o4530]='o0000;
mem_cp['o4531]='o0000;
mem_cp['o4532]='o0000;
mem_cp['o4533]='o0000;
mem_cp['o4534]='o0000;
mem_cp['o4535]='o0000;
mem_cp['o4536]='o0000;
mem_cp['o4537]='o0000;
mem_cp['o4540]='o0000;
mem_cp['o4541]='o0000;
mem_cp['o4542]='o0000;
mem_cp['o4543]='o0000;
mem_cp['o4544]='o0000;
mem_cp['o4545]='o0000;
mem_cp['o4546]='o0000;
mem_cp['o4547]='o0000;
mem_cp['o4550]='o0000;
mem_cp['o4551]='o0000;
mem_cp['o4552]='o0000;
mem_cp['o4553]='o0000;
mem_cp['o4554]='o0000;
mem_cp['o4555]='o0000;
mem_cp['o4556]='o0000;
mem_cp['o4557]='o0000;
mem_cp['o4560]='o0000;
mem_cp['o4561]='o0000;
mem_cp['o4562]='o0000;
mem_cp['o4563]='o0000;
mem_cp['o4564]='o0000;
mem_cp['o4565]='o0000;
mem_cp['o4566]='o0000;
mem_cp['o4567]='o0000;
mem_cp['o4570]='o0000;
mem_cp['o4571]='o0000;
mem_cp['o4572]='o0000;
mem_cp['o4573]='o0000;
mem_cp['o4574]='o0000;
mem_cp['o4575]='o0000;
mem_cp['o4576]='o0000;
mem_cp['o4577]='o0000;
mem_cp['o4600]='o0000;
mem_cp['o4601]='o0000;
mem_cp['o4602]='o0000;
mem_cp['o4603]='o0000;
mem_cp['o4604]='o0000;
mem_cp['o4605]='o0000;
mem_cp['o4606]='o0000;
mem_cp['o4607]='o0000;
mem_cp['o4610]='o0000;
mem_cp['o4611]='o0000;
mem_cp['o4612]='o0000;
mem_cp['o4613]='o0000;
mem_cp['o4614]='o0000;
mem_cp['o4615]='o0000;
mem_cp['o4616]='o0000;
mem_cp['o4617]='o0000;
mem_cp['o4620]='o0000;
mem_cp['o4621]='o0000;
mem_cp['o4622]='o0000;
mem_cp['o4623]='o0000;
mem_cp['o4624]='o0000;
mem_cp['o4625]='o0000;
mem_cp['o4626]='o0000;
mem_cp['o4627]='o0000;
mem_cp['o4630]='o0000;
mem_cp['o4631]='o0000;
mem_cp['o4632]='o0000;
mem_cp['o4633]='o0000;
mem_cp['o4634]='o0000;
mem_cp['o4635]='o0000;
mem_cp['o4636]='o0000;
mem_cp['o4637]='o0000;
mem_cp['o4640]='o0000;
mem_cp['o4641]='o0000;
mem_cp['o4642]='o0000;
mem_cp['o4643]='o0000;
mem_cp['o4644]='o0000;
mem_cp['o4645]='o0000;
mem_cp['o4646]='o0000;
mem_cp['o4647]='o0000;
mem_cp['o4650]='o0000;
mem_cp['o4651]='o0000;
mem_cp['o4652]='o0000;
mem_cp['o4653]='o0000;
mem_cp['o4654]='o0000;
mem_cp['o4655]='o0000;
mem_cp['o4656]='o0000;
mem_cp['o4657]='o0000;
mem_cp['o4660]='o0000;
mem_cp['o4661]='o0000;
mem_cp['o4662]='o0000;
mem_cp['o4663]='o0000;
mem_cp['o4664]='o0000;
mem_cp['o4665]='o0000;
mem_cp['o4666]='o0000;
mem_cp['o4667]='o0000;
mem_cp['o4670]='o0000;
mem_cp['o4671]='o0000;
mem_cp['o4672]='o0000;
mem_cp['o4673]='o0000;
mem_cp['o4674]='o0000;
mem_cp['o4675]='o0000;
mem_cp['o4676]='o0000;
mem_cp['o4677]='o0000;
mem_cp['o4700]='o0000;
mem_cp['o4701]='o0000;
mem_cp['o4702]='o0000;
mem_cp['o4703]='o0000;
mem_cp['o4704]='o0000;
mem_cp['o4705]='o0000;
mem_cp['o4706]='o0000;
mem_cp['o4707]='o0000;
mem_cp['o4710]='o0000;
mem_cp['o4711]='o0000;
mem_cp['o4712]='o0000;
mem_cp['o4713]='o0000;
mem_cp['o4714]='o0000;
mem_cp['o4715]='o0000;
mem_cp['o4716]='o0000;
mem_cp['o4717]='o0000;
mem_cp['o4720]='o0000;
mem_cp['o4721]='o0000;
mem_cp['o4722]='o0000;
mem_cp['o4723]='o0000;
mem_cp['o4724]='o0000;
mem_cp['o4725]='o0000;
mem_cp['o4726]='o0000;
mem_cp['o4727]='o0000;
mem_cp['o4730]='o0000;
mem_cp['o4731]='o0000;
mem_cp['o4732]='o0000;
mem_cp['o4733]='o0000;
mem_cp['o4734]='o0000;
mem_cp['o4735]='o0000;
mem_cp['o4736]='o0000;
mem_cp['o4737]='o0000;
mem_cp['o4740]='o0000;
mem_cp['o4741]='o0000;
mem_cp['o4742]='o0000;
mem_cp['o4743]='o0000;
mem_cp['o4744]='o0000;
mem_cp['o4745]='o0000;
mem_cp['o4746]='o0000;
mem_cp['o4747]='o0000;
mem_cp['o4750]='o0000;
mem_cp['o4751]='o0000;
mem_cp['o4752]='o0000;
mem_cp['o4753]='o0000;
mem_cp['o4754]='o0000;
mem_cp['o4755]='o0000;
mem_cp['o4756]='o0000;
mem_cp['o4757]='o0000;
mem_cp['o4760]='o0000;
mem_cp['o4761]='o0000;
mem_cp['o4762]='o0000;
mem_cp['o4763]='o0000;
mem_cp['o4764]='o0000;
mem_cp['o4765]='o0000;
mem_cp['o4766]='o0000;
mem_cp['o4767]='o0000;
mem_cp['o4770]='o0000;
mem_cp['o4771]='o0000;
mem_cp['o4772]='o0000;
mem_cp['o4773]='o0000;
mem_cp['o4774]='o0000;
mem_cp['o4775]='o0000;
mem_cp['o4776]='o0000;
mem_cp['o4777]='o0000;
mem_cp['o5000]='o3001;
mem_cp['o5001]='o6004;
mem_cp['o5002]='o0316;
mem_cp['o5003]='o3002;
mem_cp['o5004]='o7100;
mem_cp['o5005]='o6214;
mem_cp['o5006]='o7010;
mem_cp['o5007]='o7012;
mem_cp['o5010]='o6224;
mem_cp['o5011]='o1002;
mem_cp['o5012]='o3002;
mem_cp['o5013]='o6224;
mem_cp['o5014]='o1317;
mem_cp['o5015]='o3216;
mem_cp['o5016]='o7000;
mem_cp['o5017]='o4720;
mem_cp['o5020]='o7200;
mem_cp['o5021]='o1321;
mem_cp['o5022]='o3140;
mem_cp['o5023]='o1321;
mem_cp['o5024]='o3142;
mem_cp['o5025]='o1321;
mem_cp['o5026]='o3143;
mem_cp['o5027]='o1322;
mem_cp['o5030]='o3017;
mem_cp['o5031]='o4503;
mem_cp['o5032]='o6224;
mem_cp['o5033]='o7012;
mem_cp['o5034]='o7010;
mem_cp['o5035]='o1323;
mem_cp['o5036]='o3144;
mem_cp['o5037]='o4502;
mem_cp['o5040]='o7200;
mem_cp['o5041]='o1000;
mem_cp['o5042]='o3146;
mem_cp['o5043]='o4514;
mem_cp['o5044]='o4515;
mem_cp['o5045]='o5724;
mem_cp['o5046]='o7200;
mem_cp['o5047]='o1325;
mem_cp['o5050]='o3017;
mem_cp['o5051]='o4503;
mem_cp['o5052]='o4513;
mem_cp['o5053]='o7200;
mem_cp['o5054]='o1326;
mem_cp['o5055]='o3017;
mem_cp['o5056]='o4510;
mem_cp['o5057]='o4511;
mem_cp['o5060]='o7200;
mem_cp['o5061]='o1144;
mem_cp['o5062]='o7450;
mem_cp['o5063]='o5246;
mem_cp['o5064]='o1327;
mem_cp['o5065]='o7450;
mem_cp['o5066]='o5730;
mem_cp['o5067]='o1331;
mem_cp['o5070]='o7450;
mem_cp['o5071]='o5732;
mem_cp['o5072]='o1333;
mem_cp['o5073]='o7450;
mem_cp['o5074]='o5734;
mem_cp['o5075]='o1335;
mem_cp['o5076]='o7450;
mem_cp['o5077]='o5736;
mem_cp['o5100]='o1337;
mem_cp['o5101]='o7450;
mem_cp['o5102]='o5740;
mem_cp['o5103]='o1341;
mem_cp['o5104]='o7450;
mem_cp['o5105]='o5742;
mem_cp['o5106]='o1333;
mem_cp['o5107]='o7450;
mem_cp['o5110]='o5743;
mem_cp['o5111]='o7200;
mem_cp['o5112]='o1344;
mem_cp['o5113]='o3017;
mem_cp['o5114]='o4503;
mem_cp['o5115]='o5246;
mem_cp['o5116]='o7700;
mem_cp['o5117]='o6201;
mem_cp['o5120]='o7400;
mem_cp['o5121]='o0000;
mem_cp['o5122]='o7224;
mem_cp['o5123]='o0060;
mem_cp['o5124]='o5216;
mem_cp['o5125]='o7301;
mem_cp['o5126]='o0117;
mem_cp['o5127]='o7674;
mem_cp['o5130]='o5400;
mem_cp['o5131]='o7775;
mem_cp['o5132]='o6000;
mem_cp['o5133]='o7764;
mem_cp['o5134]='o6040;
mem_cp['o5135]='o0007;
mem_cp['o5136]='o6400;
mem_cp['o5137]='o7765;
mem_cp['o5140]='o5275;
mem_cp['o5141]='o0021;
mem_cp['o5142]='o5247;
mem_cp['o5143]='o5200;
mem_cp['o5144]='o7321;
mem_cp['o5145]='o0000;
mem_cp['o5146]='o0000;
mem_cp['o5147]='o0000;
mem_cp['o5150]='o0000;
mem_cp['o5151]='o0000;
mem_cp['o5152]='o0000;
mem_cp['o5153]='o0000;
mem_cp['o5154]='o0000;
mem_cp['o5155]='o0000;
mem_cp['o5156]='o0000;
mem_cp['o5157]='o0000;
mem_cp['o5160]='o0000;
mem_cp['o5161]='o0000;
mem_cp['o5162]='o0000;
mem_cp['o5163]='o0000;
mem_cp['o5164]='o0000;
mem_cp['o5165]='o0000;
mem_cp['o5166]='o0000;
mem_cp['o5167]='o0000;
mem_cp['o5170]='o0000;
mem_cp['o5171]='o0000;
mem_cp['o5172]='o0000;
mem_cp['o5173]='o0000;
mem_cp['o5174]='o0000;
mem_cp['o5175]='o0000;
mem_cp['o5176]='o0000;
mem_cp['o5177]='o0000;
mem_cp['o5200]='o2017;
mem_cp['o5201]='o4510;
mem_cp['o5202]='o4512;
mem_cp['o5203]='o4510;
mem_cp['o5204]='o7200;
mem_cp['o5205]='o1144;
mem_cp['o5206]='o7440;
mem_cp['o5207]='o5507;
mem_cp['o5210]='o1145;
mem_cp['o5211]='o7450;
mem_cp['o5212]='o5216;
mem_cp['o5213]='o7200;
mem_cp['o5214]='o1146;
mem_cp['o5215]='o3001;
mem_cp['o5216]='o7200;
mem_cp['o5217]='o1314;
mem_cp['o5220]='o3017;
mem_cp['o5221]='o4503;
mem_cp['o5222]='o7200;
mem_cp['o5223]='o1001;
mem_cp['o5224]='o3146;
mem_cp['o5225]='o4514;
mem_cp['o5226]='o1315;
mem_cp['o5227]='o3017;
mem_cp['o5230]='o4503;
mem_cp['o5231]='o7200;
mem_cp['o5232]='o1002;
mem_cp['o5233]='o3146;
mem_cp['o5234]='o4514;
mem_cp['o5235]='o1316;
mem_cp['o5236]='o3017;
mem_cp['o5237]='o4503;
mem_cp['o5240]='o7200;
mem_cp['o5241]='o7404;
mem_cp['o5242]='o3146;
mem_cp['o5243]='o4514;
mem_cp['o5244]='o4515;
mem_cp['o5245]='o5501;
mem_cp['o5246]='o5501;
mem_cp['o5247]='o2017;
mem_cp['o5250]='o4510;
mem_cp['o5251]='o4512;
mem_cp['o5252]='o4510;
mem_cp['o5253]='o7200;
mem_cp['o5254]='o1144;
mem_cp['o5255]='o7440;
mem_cp['o5256]='o5507;
mem_cp['o5257]='o1145;
mem_cp['o5260]='o7450;
mem_cp['o5261]='o5274;
mem_cp['o5262]='o7300;
mem_cp['o5263]='o1146;
mem_cp['o5264]='o3002;
mem_cp['o5265]='o1002;
mem_cp['o5266]='o7004;
mem_cp['o5267]='o7006;
mem_cp['o5270]='o0317;
mem_cp['o5271]='o1320;
mem_cp['o5272]='o3273;
mem_cp['o5273]='o7000;
mem_cp['o5274]='o5216;
mem_cp['o5275]='o2017;
mem_cp['o5276]='o4510;
mem_cp['o5277]='o4512;
mem_cp['o5300]='o4510;
mem_cp['o5301]='o7200;
mem_cp['o5302]='o1144;
mem_cp['o5303]='o7440;
mem_cp['o5304]='o5507;
mem_cp['o5305]='o1145;
mem_cp['o5306]='o7450;
mem_cp['o5307]='o5313;
mem_cp['o5310]='o7200;
mem_cp['o5311]='o1146;
mem_cp['o5312]='o6301;
mem_cp['o5313]='o5216;
mem_cp['o5314]='o7345;
mem_cp['o5315]='o7351;
mem_cp['o5316]='o7365;
mem_cp['o5317]='o0070;
mem_cp['o5320]='o6201;
mem_cp['o5321]='o0000;
mem_cp['o5322]='o0000;
mem_cp['o5323]='o0000;
mem_cp['o5324]='o0000;
mem_cp['o5325]='o0000;
mem_cp['o5326]='o0000;
mem_cp['o5327]='o0000;
mem_cp['o5330]='o0000;
mem_cp['o5331]='o0000;
mem_cp['o5332]='o0000;
mem_cp['o5333]='o0000;
mem_cp['o5334]='o0000;
mem_cp['o5335]='o0000;
mem_cp['o5336]='o0000;
mem_cp['o5337]='o0000;
mem_cp['o5340]='o0000;
mem_cp['o5341]='o0000;
mem_cp['o5342]='o0000;
mem_cp['o5343]='o0000;
mem_cp['o5344]='o0000;
mem_cp['o5345]='o0000;
mem_cp['o5346]='o0000;
mem_cp['o5347]='o0000;
mem_cp['o5350]='o0000;
mem_cp['o5351]='o0000;
mem_cp['o5352]='o0000;
mem_cp['o5353]='o0000;
mem_cp['o5354]='o0000;
mem_cp['o5355]='o0000;
mem_cp['o5356]='o0000;
mem_cp['o5357]='o0000;
mem_cp['o5360]='o0000;
mem_cp['o5361]='o0000;
mem_cp['o5362]='o0000;
mem_cp['o5363]='o0000;
mem_cp['o5364]='o0000;
mem_cp['o5365]='o0000;
mem_cp['o5366]='o0000;
mem_cp['o5367]='o0000;
mem_cp['o5370]='o0000;
mem_cp['o5371]='o0000;
mem_cp['o5372]='o0000;
mem_cp['o5373]='o0000;
mem_cp['o5374]='o0000;
mem_cp['o5375]='o0000;
mem_cp['o5376]='o0000;
mem_cp['o5377]='o0000;
mem_cp['o5400]='o2017;
mem_cp['o5401]='o4510;
mem_cp['o5402]='o4512;
mem_cp['o5403]='o7200;
mem_cp['o5404]='o1145;
mem_cp['o5405]='o7440;
mem_cp['o5406]='o5220;
mem_cp['o5407]='o4510;
mem_cp['o5410]='o7200;
mem_cp['o5411]='o1144;
mem_cp['o5412]='o7440;
mem_cp['o5413]='o5507;
mem_cp['o5414]='o1140;
mem_cp['o5415]='o1332;
mem_cp['o5416]='o3141;
mem_cp['o5417]='o5260;
mem_cp['o5420]='o7200;
mem_cp['o5421]='o1146;
mem_cp['o5422]='o3140;
mem_cp['o5423]='o4510;
mem_cp['o5424]='o7200;
mem_cp['o5425]='o1144;
mem_cp['o5426]='o1333;
mem_cp['o5427]='o7450;
mem_cp['o5430]='o5241;
mem_cp['o5431]='o1334;
mem_cp['o5432]='o7440;
mem_cp['o5433]='o5507;
mem_cp['o5434]='o7200;
mem_cp['o5435]='o1140;
mem_cp['o5436]='o1332;
mem_cp['o5437]='o3141;
mem_cp['o5440]='o5260;
mem_cp['o5441]='o2017;
mem_cp['o5442]='o4510;
mem_cp['o5443]='o4512;
mem_cp['o5444]='o4510;
mem_cp['o5445]='o7200;
mem_cp['o5446]='o1145;
mem_cp['o5447]='o7450;
mem_cp['o5450]='o5507;
mem_cp['o5451]='o7200;
mem_cp['o5452]='o1144;
mem_cp['o5453]='o7440;
mem_cp['o5454]='o5507;
mem_cp['o5455]='o7001;
mem_cp['o5456]='o1146;
mem_cp['o5457]='o3141;
mem_cp['o5460]='o7200;
mem_cp['o5461]='o1140;
mem_cp['o5462]='o0335;
mem_cp['o5463]='o1336;
mem_cp['o5464]='o3016;
mem_cp['o5465]='o3147;
mem_cp['o5466]='o4311;
mem_cp['o5467]='o4505;
mem_cp['o5470]='o7200;
mem_cp['o5471]='o1144;
mem_cp['o5472]='o7440;
mem_cp['o5473]='o5304;
mem_cp['o5474]='o1147;
mem_cp['o5475]='o1337;
mem_cp['o5476]='o7510;
mem_cp['o5477]='o5266;
mem_cp['o5500]='o7200;
mem_cp['o5501]='o1141;
mem_cp['o5502]='o3140;
mem_cp['o5503]='o5501;
mem_cp['o5504]='o7200;
mem_cp['o5505]='o1016;
mem_cp['o5506]='o3140;
mem_cp['o5507]='o4504;
mem_cp['o5510]='o5501;
mem_cp['o5511]='o0000;
mem_cp['o5512]='o7200;
mem_cp['o5513]='o1016;
mem_cp['o5514]='o7001;
mem_cp['o5515]='o3146;
mem_cp['o5516]='o4514;
mem_cp['o5517]='o1340;
mem_cp['o5520]='o3017;
mem_cp['o5521]='o4503;
mem_cp['o5522]='o7200;
mem_cp['o5523]='o1335;
mem_cp['o5524]='o3145;
mem_cp['o5525]='o4741;
mem_cp['o5526]='o2145;
mem_cp['o5527]='o5325;
mem_cp['o5530]='o4515;
mem_cp['o5531]='o5711;
mem_cp['o5532]='o0100;
mem_cp['o5533]='o7724;
mem_cp['o5534]='o0054;
mem_cp['o5535]='o7770;
mem_cp['o5536]='o7777;
mem_cp['o5537]='o7776;
mem_cp['o5540]='o7331;
mem_cp['o5541]='o5600;
mem_cp['o5542]='o0000;
mem_cp['o5543]='o0000;
mem_cp['o5544]='o0000;
mem_cp['o5545]='o0000;
mem_cp['o5546]='o0000;
mem_cp['o5547]='o0000;
mem_cp['o5550]='o0000;
mem_cp['o5551]='o0000;
mem_cp['o5552]='o0000;
mem_cp['o5553]='o0000;
mem_cp['o5554]='o0000;
mem_cp['o5555]='o0000;
mem_cp['o5556]='o0000;
mem_cp['o5557]='o0000;
mem_cp['o5560]='o0000;
mem_cp['o5561]='o0000;
mem_cp['o5562]='o0000;
mem_cp['o5563]='o0000;
mem_cp['o5564]='o0000;
mem_cp['o5565]='o0000;
mem_cp['o5566]='o0000;
mem_cp['o5567]='o0000;
mem_cp['o5570]='o0000;
mem_cp['o5571]='o0000;
mem_cp['o5572]='o0000;
mem_cp['o5573]='o0000;
mem_cp['o5574]='o0000;
mem_cp['o5575]='o0000;
mem_cp['o5576]='o0000;
mem_cp['o5577]='o0000;
mem_cp['o5600]='o0000;
mem_cp['o5601]='o7200;
mem_cp['o5602]='o1246;
mem_cp['o5603]='o3144;
mem_cp['o5604]='o4502;
mem_cp['o5605]='o7200;
mem_cp['o5606]='o1147;
mem_cp['o5607]='o7440;
mem_cp['o5610]='o5230;
mem_cp['o5611]='o1016;
mem_cp['o5612]='o7040;
mem_cp['o5613]='o1140;
mem_cp['o5614]='o7450;
mem_cp['o5615]='o5227;
mem_cp['o5616]='o7200;
mem_cp['o5617]='o1247;
mem_cp['o5620]='o3017;
mem_cp['o5621]='o4503;
mem_cp['o5622]='o7200;
mem_cp['o5623]='o1016;
mem_cp['o5624]='o7001;
mem_cp['o5625]='o3016;
mem_cp['o5626]='o5600;
mem_cp['o5627]='o2147;
mem_cp['o5630]='o7240;
mem_cp['o5631]='o1147;
mem_cp['o5632]='o7440;
mem_cp['o5633]='o5216;
mem_cp['o5634]='o7200;
mem_cp['o5635]='o1416;
mem_cp['o5636]='o3146;
mem_cp['o5637]='o4514;
mem_cp['o5640]='o1016;
mem_cp['o5641]='o7040;
mem_cp['o5642]='o1141;
mem_cp['o5643]='o7450;
mem_cp['o5644]='o2147;
mem_cp['o5645]='o5600;
mem_cp['o5646]='o0040;
mem_cp['o5647]='o7340;
mem_cp['o5650]='o0000;
mem_cp['o5651]='o0000;
mem_cp['o5652]='o0000;
mem_cp['o5653]='o0000;
mem_cp['o5654]='o0000;
mem_cp['o5655]='o0000;
mem_cp['o5656]='o0000;
mem_cp['o5657]='o0000;
mem_cp['o5660]='o0000;
mem_cp['o5661]='o0000;
mem_cp['o5662]='o0000;
mem_cp['o5663]='o0000;
mem_cp['o5664]='o0000;
mem_cp['o5665]='o0000;
mem_cp['o5666]='o0000;
mem_cp['o5667]='o0000;
mem_cp['o5670]='o0000;
mem_cp['o5671]='o0000;
mem_cp['o5672]='o0000;
mem_cp['o5673]='o0000;
mem_cp['o5674]='o0000;
mem_cp['o5675]='o0000;
mem_cp['o5676]='o0000;
mem_cp['o5677]='o0000;
mem_cp['o5700]='o0000;
mem_cp['o5701]='o0000;
mem_cp['o5702]='o0000;
mem_cp['o5703]='o0000;
mem_cp['o5704]='o0000;
mem_cp['o5705]='o0000;
mem_cp['o5706]='o0000;
mem_cp['o5707]='o0000;
mem_cp['o5710]='o0000;
mem_cp['o5711]='o0000;
mem_cp['o5712]='o0000;
mem_cp['o5713]='o0000;
mem_cp['o5714]='o0000;
mem_cp['o5715]='o0000;
mem_cp['o5716]='o0000;
mem_cp['o5717]='o0000;
mem_cp['o5720]='o0000;
mem_cp['o5721]='o0000;
mem_cp['o5722]='o0000;
mem_cp['o5723]='o0000;
mem_cp['o5724]='o0000;
mem_cp['o5725]='o0000;
mem_cp['o5726]='o0000;
mem_cp['o5727]='o0000;
mem_cp['o5730]='o0000;
mem_cp['o5731]='o0000;
mem_cp['o5732]='o0000;
mem_cp['o5733]='o0000;
mem_cp['o5734]='o0000;
mem_cp['o5735]='o0000;
mem_cp['o5736]='o0000;
mem_cp['o5737]='o0000;
mem_cp['o5740]='o0000;
mem_cp['o5741]='o0000;
mem_cp['o5742]='o0000;
mem_cp['o5743]='o0000;
mem_cp['o5744]='o0000;
mem_cp['o5745]='o0000;
mem_cp['o5746]='o0000;
mem_cp['o5747]='o0000;
mem_cp['o5750]='o0000;
mem_cp['o5751]='o0000;
mem_cp['o5752]='o0000;
mem_cp['o5753]='o0000;
mem_cp['o5754]='o0000;
mem_cp['o5755]='o0000;
mem_cp['o5756]='o0000;
mem_cp['o5757]='o0000;
mem_cp['o5760]='o0000;
mem_cp['o5761]='o0000;
mem_cp['o5762]='o0000;
mem_cp['o5763]='o0000;
mem_cp['o5764]='o0000;
mem_cp['o5765]='o0000;
mem_cp['o5766]='o0000;
mem_cp['o5767]='o0000;
mem_cp['o5770]='o0000;
mem_cp['o5771]='o0000;
mem_cp['o5772]='o0000;
mem_cp['o5773]='o0000;
mem_cp['o5774]='o0000;
mem_cp['o5775]='o0000;
mem_cp['o5776]='o0000;
mem_cp['o5777]='o0000;
mem_cp['o6000]='o2017;
mem_cp['o6001]='o4510;
mem_cp['o6002]='o4512;
mem_cp['o6003]='o4510;
mem_cp['o6004]='o7200;
mem_cp['o6005]='o1144;
mem_cp['o6006]='o7440;
mem_cp['o6007]='o5507;
mem_cp['o6010]='o1145;
mem_cp['o6011]='o7450;
mem_cp['o6012]='o5216;
mem_cp['o6013]='o7200;
mem_cp['o6014]='o1146;
mem_cp['o6015]='o3000;
mem_cp['o6016]='o1002;
mem_cp['o6017]='o7004;
mem_cp['o6020]='o7006;
mem_cp['o6021]='o0340;
mem_cp['o6022]='o1341;
mem_cp['o6023]='o3224;
mem_cp['o6024]='o7000;
mem_cp['o6025]='o1002;
mem_cp['o6026]='o7004;
mem_cp['o6027]='o1002;
mem_cp['o6030]='o0340;
mem_cp['o6031]='o1342;
mem_cp['o6032]='o3233;
mem_cp['o6033]='o7000;
mem_cp['o6034]='o7200;
mem_cp['o6035]='o1001;
mem_cp['o6036]='o6001;
mem_cp['o6037]='o5400;
mem_cp['o6040]='o2017;
mem_cp['o6041]='o4510;
mem_cp['o6042]='o4512;
mem_cp['o6043]='o4510;
mem_cp['o6044]='o7200;
mem_cp['o6045]='o1144;
mem_cp['o6046]='o7440;
mem_cp['o6047]='o5507;
mem_cp['o6050]='o1145;
mem_cp['o6051]='o7450;
mem_cp['o6052]='o5256;
mem_cp['o6053]='o7200;
mem_cp['o6054]='o1146;
mem_cp['o6055]='o3142;
mem_cp['o6056]='o7200;
mem_cp['o6057]='o1142;
mem_cp['o6060]='o3146;
mem_cp['o6061]='o4514;
mem_cp['o6062]='o7200;
mem_cp['o6063]='o1343;
mem_cp['o6064]='o3017;
mem_cp['o6065]='o4503;
mem_cp['o6066]='o7200;
mem_cp['o6067]='o1542;
mem_cp['o6070]='o3146;
mem_cp['o6071]='o4514;
mem_cp['o6072]='o7200;
mem_cp['o6073]='o1344;
mem_cp['o6074]='o3144;
mem_cp['o6075]='o4502;
mem_cp['o6076]='o4513;
mem_cp['o6077]='o7200;
mem_cp['o6100]='o1345;
mem_cp['o6101]='o3017;
mem_cp['o6102]='o4510;
mem_cp['o6103]='o7200;
mem_cp['o6104]='o1144;
mem_cp['o6105]='o7440;
mem_cp['o6106]='o5312;
mem_cp['o6107]='o2142;
mem_cp['o6110]='o7000;
mem_cp['o6111]='o5256;
mem_cp['o6112]='o1346;
mem_cp['o6113]='o7440;
mem_cp['o6114]='o5321;
mem_cp['o6115]='o7240;
mem_cp['o6116]='o1142;
mem_cp['o6117]='o3142;
mem_cp['o6120]='o5256;
mem_cp['o6121]='o1347;
mem_cp['o6122]='o7440;
mem_cp['o6123]='o5325;
mem_cp['o6124]='o5501;
mem_cp['o6125]='o4512;
mem_cp['o6126]='o7200;
mem_cp['o6127]='o1145;
mem_cp['o6130]='o7450;
mem_cp['o6131]='o5507;
mem_cp['o6132]='o7200;
mem_cp['o6133]='o1146;
mem_cp['o6134]='o3542;
mem_cp['o6135]='o2142;
mem_cp['o6136]='o7000;
mem_cp['o6137]='o5256;
mem_cp['o6140]='o0070;
mem_cp['o6141]='o6201;
mem_cp['o6142]='o6202;
mem_cp['o6143]='o7334;
mem_cp['o6144]='o0040;
mem_cp['o6145]='o0117;
mem_cp['o6146]='o7723;
mem_cp['o6147]='o7777;
mem_cp['o6150]='o0000;
mem_cp['o6151]='o0000;
mem_cp['o6152]='o0000;
mem_cp['o6153]='o0000;
mem_cp['o6154]='o0000;
mem_cp['o6155]='o0000;
mem_cp['o6156]='o0000;
mem_cp['o6157]='o0000;
mem_cp['o6160]='o0000;
mem_cp['o6161]='o0000;
mem_cp['o6162]='o0000;
mem_cp['o6163]='o0000;
mem_cp['o6164]='o0000;
mem_cp['o6165]='o0000;
mem_cp['o6166]='o0000;
mem_cp['o6167]='o0000;
mem_cp['o6170]='o0000;
mem_cp['o6171]='o0000;
mem_cp['o6172]='o0000;
mem_cp['o6173]='o0000;
mem_cp['o6174]='o0000;
mem_cp['o6175]='o0000;
mem_cp['o6176]='o0000;
mem_cp['o6177]='o0000;
mem_cp['o6200]='o0000;
mem_cp['o6201]='o7200;
mem_cp['o6202]='o3146;
mem_cp['o6203]='o4213;
mem_cp['o6204]='o7200;
mem_cp['o6205]='o1146;
mem_cp['o6206]='o7106;
mem_cp['o6207]='o7106;
mem_cp['o6210]='o3146;
mem_cp['o6211]='o4213;
mem_cp['o6212]='o5600;
mem_cp['o6213]='o0000;
mem_cp['o6214]='o4504;
mem_cp['o6215]='o4511;
mem_cp['o6216]='o7200;
mem_cp['o6217]='o1144;
mem_cp['o6220]='o1246;
mem_cp['o6221]='o7510;
mem_cp['o6222]='o5245;
mem_cp['o6223]='o1247;
mem_cp['o6224]='o7510;
mem_cp['o6225]='o5240;
mem_cp['o6226]='o1250;
mem_cp['o6227]='o7510;
mem_cp['o6230]='o5245;
mem_cp['o6231]='o1251;
mem_cp['o6232]='o7500;
mem_cp['o6233]='o5245;
mem_cp['o6234]='o7200;
mem_cp['o6235]='o1144;
mem_cp['o6236]='o1252;
mem_cp['o6237]='o5243;
mem_cp['o6240]='o7200;
mem_cp['o6241]='o1144;
mem_cp['o6242]='o1246;
mem_cp['o6243]='o1146;
mem_cp['o6244]='o3146;
mem_cp['o6245]='o5613;
mem_cp['o6246]='o7720;
mem_cp['o6247]='o7766;
mem_cp['o6250]='o7771;
mem_cp['o6251]='o7772;
mem_cp['o6252]='o7711;
mem_cp['o6253]='o0000;
mem_cp['o6254]='o0000;
mem_cp['o6255]='o0000;
mem_cp['o6256]='o0000;
mem_cp['o6257]='o0000;
mem_cp['o6260]='o0000;
mem_cp['o6261]='o0000;
mem_cp['o6262]='o0000;
mem_cp['o6263]='o0000;
mem_cp['o6264]='o0000;
mem_cp['o6265]='o0000;
mem_cp['o6266]='o0000;
mem_cp['o6267]='o0000;
mem_cp['o6270]='o0000;
mem_cp['o6271]='o0000;
mem_cp['o6272]='o0000;
mem_cp['o6273]='o0000;
mem_cp['o6274]='o0000;
mem_cp['o6275]='o0000;
mem_cp['o6276]='o0000;
mem_cp['o6277]='o0000;
mem_cp['o6300]='o0000;
mem_cp['o6301]='o0000;
mem_cp['o6302]='o0000;
mem_cp['o6303]='o0000;
mem_cp['o6304]='o0000;
mem_cp['o6305]='o0000;
mem_cp['o6306]='o0000;
mem_cp['o6307]='o0000;
mem_cp['o6310]='o0000;
mem_cp['o6311]='o0000;
mem_cp['o6312]='o0000;
mem_cp['o6313]='o0000;
mem_cp['o6314]='o0000;
mem_cp['o6315]='o0000;
mem_cp['o6316]='o0000;
mem_cp['o6317]='o0000;
mem_cp['o6320]='o0000;
mem_cp['o6321]='o0000;
mem_cp['o6322]='o0000;
mem_cp['o6323]='o0000;
mem_cp['o6324]='o0000;
mem_cp['o6325]='o0000;
mem_cp['o6326]='o0000;
mem_cp['o6327]='o0000;
mem_cp['o6330]='o0000;
mem_cp['o6331]='o0000;
mem_cp['o6332]='o0000;
mem_cp['o6333]='o0000;
mem_cp['o6334]='o0000;
mem_cp['o6335]='o0000;
mem_cp['o6336]='o0000;
mem_cp['o6337]='o0000;
mem_cp['o6340]='o0000;
mem_cp['o6341]='o0000;
mem_cp['o6342]='o0000;
mem_cp['o6343]='o0000;
mem_cp['o6344]='o0000;
mem_cp['o6345]='o0000;
mem_cp['o6346]='o0000;
mem_cp['o6347]='o0000;
mem_cp['o6350]='o0000;
mem_cp['o6351]='o0000;
mem_cp['o6352]='o0000;
mem_cp['o6353]='o0000;
mem_cp['o6354]='o0000;
mem_cp['o6355]='o0000;
mem_cp['o6356]='o0000;
mem_cp['o6357]='o0000;
mem_cp['o6360]='o0000;
mem_cp['o6361]='o0000;
mem_cp['o6362]='o0000;
mem_cp['o6363]='o0000;
mem_cp['o6364]='o0000;
mem_cp['o6365]='o0000;
mem_cp['o6366]='o0000;
mem_cp['o6367]='o0000;
mem_cp['o6370]='o0000;
mem_cp['o6371]='o0000;
mem_cp['o6372]='o0000;
mem_cp['o6373]='o0000;
mem_cp['o6374]='o0000;
mem_cp['o6375]='o0000;
mem_cp['o6376]='o0000;
mem_cp['o6377]='o0000;
mem_cp['o6400]='o2017;
mem_cp['o6401]='o4510;
mem_cp['o6402]='o4512;
mem_cp['o6403]='o4510;
mem_cp['o6404]='o7200;
mem_cp['o6405]='o1144;
mem_cp['o6406]='o7440;
mem_cp['o6407]='o5507;
mem_cp['o6410]='o7240;
mem_cp['o6411]='o1146;
mem_cp['o6412]='o3016;
mem_cp['o6413]='o4504;
mem_cp['o6414]='o4511;
mem_cp['o6415]='o7200;
mem_cp['o6416]='o1144;
mem_cp['o6417]='o1367;
mem_cp['o6420]='o7450;
mem_cp['o6421]='o5234;
mem_cp['o6422]='o7200;
mem_cp['o6423]='o1144;
mem_cp['o6424]='o1370;
mem_cp['o6425]='o7450;
mem_cp['o6426]='o5213;
mem_cp['o6427]='o1371;
mem_cp['o6430]='o7450;
mem_cp['o6431]='o5213;
mem_cp['o6432]='o4504;
mem_cp['o6433]='o5222;
mem_cp['o6434]='o4772;
mem_cp['o6435]='o7200;
mem_cp['o6436]='o1146;
mem_cp['o6437]='o3150;
mem_cp['o6440]='o1146;
mem_cp['o6441]='o7110;
mem_cp['o6442]='o7430;
mem_cp['o6443]='o5362;
mem_cp['o6444]='o7041;
mem_cp['o6445]='o3145;
mem_cp['o6446]='o4772;
mem_cp['o6447]='o7200;
mem_cp['o6450]='o1146;
mem_cp['o6451]='o1150;
mem_cp['o6452]='o3150;
mem_cp['o6453]='o1146;
mem_cp['o6454]='o7002;
mem_cp['o6455]='o7104;
mem_cp['o6456]='o0373;
mem_cp['o6457]='o3017;
mem_cp['o6460]='o4772;
mem_cp['o6461]='o7200;
mem_cp['o6462]='o1146;
mem_cp['o6463]='o1150;
mem_cp['o6464]='o3150;
mem_cp['o6465]='o1146;
mem_cp['o6466]='o7110;
mem_cp['o6467]='o7430;
mem_cp['o6470]='o5507;
mem_cp['o6471]='o1017;
mem_cp['o6472]='o1016;
mem_cp['o6473]='o3017;
mem_cp['o6474]='o4772;
mem_cp['o6475]='o7200;
mem_cp['o6476]='o1146;
mem_cp['o6477]='o1150;
mem_cp['o6500]='o3150;
mem_cp['o6501]='o7040;
mem_cp['o6502]='o1146;
mem_cp['o6503]='o7450;
mem_cp['o6504]='o5311;
mem_cp['o6505]='o7001;
mem_cp['o6506]='o7450;
mem_cp['o6507]='o5311;
mem_cp['o6510]='o5232;
mem_cp['o6511]='o1146;
mem_cp['o6512]='o3147;
mem_cp['o6513]='o1145;
mem_cp['o6514]='o7450;
mem_cp['o6515]='o5345;
mem_cp['o6516]='o4772;
mem_cp['o6517]='o7200;
mem_cp['o6520]='o1146;
mem_cp['o6521]='o1150;
mem_cp['o6522]='o3150;
mem_cp['o6523]='o1146;
mem_cp['o6524]='o7002;
mem_cp['o6525]='o7006;
mem_cp['o6526]='o0373;
mem_cp['o6527]='o3120;
mem_cp['o6530]='o4772;
mem_cp['o6531]='o7200;
mem_cp['o6532]='o1146;
mem_cp['o6533]='o1150;
mem_cp['o6534]='o3150;
mem_cp['o6535]='o1147;
mem_cp['o6536]='o7440;
mem_cp['o6537]='o5343;
mem_cp['o6540]='o1146;
mem_cp['o6541]='o1120;
mem_cp['o6542]='o3417;
mem_cp['o6543]='o2145;
mem_cp['o6544]='o5316;
mem_cp['o6545]='o4772;
mem_cp['o6546]='o7200;
mem_cp['o6547]='o1146;
mem_cp['o6550]='o1150;
mem_cp['o6551]='o0374;
mem_cp['o6552]='o7440;
mem_cp['o6553]='o5362;
mem_cp['o6554]='o4775;
mem_cp['o6555]='o7240;
mem_cp['o6556]='o1147;
mem_cp['o6557]='o7440;
mem_cp['o6560]='o5232;
mem_cp['o6561]='o5501;
mem_cp['o6562]='o7200;
mem_cp['o6563]='o1376;
mem_cp['o6564]='o3017;
mem_cp['o6565]='o4503;
mem_cp['o6566]='o5501;
mem_cp['o6567]='o7706;
mem_cp['o6570]='o7763;
mem_cp['o6571]='o0003;
mem_cp['o6572]='o6200;
mem_cp['o6573]='o7400;
mem_cp['o6574]='o0377;
mem_cp['o6575]='o7216;
mem_cp['o6576]='o7304;
mem_cp['o6577]='o0000;
mem_cp['o6600]='o0000;
mem_cp['o6601]='o7200;
mem_cp['o6602]='o1146;
mem_cp['o6603]='o7010;
mem_cp['o6604]='o7012;
mem_cp['o6605]='o0347;
mem_cp['o6606]='o1350;
mem_cp['o6607]='o3144;
mem_cp['o6610]='o4502;
mem_cp['o6611]='o7200;
mem_cp['o6612]='o1146;
mem_cp['o6613]='o0347;
mem_cp['o6614]='o1350;
mem_cp['o6615]='o3144;
mem_cp['o6616]='o4502;
mem_cp['o6617]='o5600;
mem_cp['o6620]='o0000;
mem_cp['o6621]='o7200;
mem_cp['o6622]='o1146;
mem_cp['o6623]='o7002;
mem_cp['o6624]='o3146;
mem_cp['o6625]='o4200;
mem_cp['o6626]='o7200;
mem_cp['o6627]='o1146;
mem_cp['o6630]='o7002;
mem_cp['o6631]='o3146;
mem_cp['o6632]='o4200;
mem_cp['o6633]='o5620;
mem_cp['o6634]='o0000;
mem_cp['o6635]='o7200;
mem_cp['o6636]='o1351;
mem_cp['o6637]='o3144;
mem_cp['o6640]='o4502;
mem_cp['o6641]='o7200;
mem_cp['o6642]='o1352;
mem_cp['o6643]='o3144;
mem_cp['o6644]='o4502;
mem_cp['o6645]='o5634;
mem_cp['o6646]='o0000;
mem_cp['o6647]='o7200;
mem_cp['o6650]='o3145;
mem_cp['o6651]='o1353;
mem_cp['o6652]='o3017;
mem_cp['o6653]='o4504;
mem_cp['o6654]='o7200;
mem_cp['o6655]='o1144;
mem_cp['o6656]='o1354;
mem_cp['o6657]='o7450;
mem_cp['o6660]='o5343;
mem_cp['o6661]='o1355;
mem_cp['o6662]='o7450;
mem_cp['o6663]='o5343;
mem_cp['o6664]='o1356;
mem_cp['o6665]='o7450;
mem_cp['o6666]='o5315;
mem_cp['o6667]='o1357;
mem_cp['o6670]='o7450;
mem_cp['o6671]='o5315;
mem_cp['o6672]='o1360;
mem_cp['o6673]='o7510;
mem_cp['o6674]='o5253;
mem_cp['o6675]='o1361;
mem_cp['o6676]='o7500;
mem_cp['o6677]='o5253;
mem_cp['o6700]='o7200;
mem_cp['o6701]='o1145;
mem_cp['o6702]='o1362;
mem_cp['o6703]='o7500;
mem_cp['o6704]='o5253;
mem_cp['o6705]='o7200;
mem_cp['o6706]='o1144;
mem_cp['o6707]='o4161;
mem_cp['o6710]='o1144;
mem_cp['o6711]='o4502;
mem_cp['o6712]='o2145;
mem_cp['o6713]='o7000;
mem_cp['o6714]='o5253;
mem_cp['o6715]='o7200;
mem_cp['o6716]='o1145;
mem_cp['o6717]='o7450;
mem_cp['o6720]='o5253;
mem_cp['o6721]='o7240;
mem_cp['o6722]='o1145;
mem_cp['o6723]='o3145;
mem_cp['o6724]='o7240;
mem_cp['o6725]='o1017;
mem_cp['o6726]='o3017;
mem_cp['o6727]='o1363;
mem_cp['o6730]='o3144;
mem_cp['o6731]='o4502;
mem_cp['o6732]='o7200;
mem_cp['o6733]='o1364;
mem_cp['o6734]='o3144;
mem_cp['o6735]='o4502;
mem_cp['o6736]='o7200;
mem_cp['o6737]='o1363;
mem_cp['o6740]='o3144;
mem_cp['o6741]='o4502;
mem_cp['o6742]='o5253;
mem_cp['o6743]='o4234;
mem_cp['o6744]='o7200;
mem_cp['o6745]='o4161;
mem_cp['o6746]='o5646;
mem_cp['o6747]='o0007;
mem_cp['o6750]='o0060;
mem_cp['o6751]='o0015;
mem_cp['o6752]='o0012;
mem_cp['o6753]='o0117;
mem_cp['o6754]='o7763;
mem_cp['o6755]='o0003;
mem_cp['o6756]='o0002;
mem_cp['o6757]='o7611;
mem_cp['o6760]='o0137;
mem_cp['o6761]='o7640;
mem_cp['o6762]='o7761;
mem_cp['o6763]='o0010;
mem_cp['o6764]='o0040;
mem_cp['o6765]='o0000;
mem_cp['o6766]='o0000;
mem_cp['o6767]='o0000;
mem_cp['o6770]='o0000;
mem_cp['o6771]='o0000;
mem_cp['o6772]='o0000;
mem_cp['o6773]='o0000;
mem_cp['o6774]='o0000;
mem_cp['o6775]='o0000;
mem_cp['o6776]='o0000;
mem_cp['o6777]='o0000;
mem_cp['o7000]='o0000;
mem_cp['o7001]='o7200;
mem_cp['o7002]='o4151;
mem_cp['o7003]='o3144;
mem_cp['o7004]='o1144;
mem_cp['o7005]='o1273;
mem_cp['o7006]='o7450;
mem_cp['o7007]='o5201;
mem_cp['o7010]='o7240;
mem_cp['o7011]='o1017;
mem_cp['o7012]='o3017;
mem_cp['o7013]='o5600;
mem_cp['o7014]='o0000;
mem_cp['o7015]='o7200;
mem_cp['o7016]='o1144;
mem_cp['o7017]='o1274;
mem_cp['o7020]='o7510;
mem_cp['o7021]='o5614;
mem_cp['o7022]='o7200;
mem_cp['o7023]='o1144;
mem_cp['o7024]='o1275;
mem_cp['o7025]='o7540;
mem_cp['o7026]='o5614;
mem_cp['o7027]='o1276;
mem_cp['o7030]='o3144;
mem_cp['o7031]='o5614;
mem_cp['o7032]='o0000;
mem_cp['o7033]='o7200;
mem_cp['o7034]='o3145;
mem_cp['o7035]='o3146;
mem_cp['o7036]='o7200;
mem_cp['o7037]='o4151;
mem_cp['o7040]='o3144;
mem_cp['o7041]='o4214;
mem_cp['o7042]='o7200;
mem_cp['o7043]='o1144;
mem_cp['o7044]='o1277;
mem_cp['o7045]='o7540;
mem_cp['o7046]='o5267;
mem_cp['o7047]='o7200;
mem_cp['o7050]='o1144;
mem_cp['o7051]='o1300;
mem_cp['o7052]='o7510;
mem_cp['o7053]='o5267;
mem_cp['o7054]='o0301;
mem_cp['o7055]='o3144;
mem_cp['o7056]='o1146;
mem_cp['o7057]='o7004;
mem_cp['o7060]='o7006;
mem_cp['o7061]='o0302;
mem_cp['o7062]='o1144;
mem_cp['o7063]='o3146;
mem_cp['o7064]='o2145;
mem_cp['o7065]='o7000;
mem_cp['o7066]='o5236;
mem_cp['o7067]='o7240;
mem_cp['o7070]='o1017;
mem_cp['o7071]='o3017;
mem_cp['o7072]='o5632;
mem_cp['o7073]='o7740;
mem_cp['o7074]='o7637;
mem_cp['o7075]='o7606;
mem_cp['o7076]='o0132;
mem_cp['o7077]='o7707;
mem_cp['o7100]='o7720;
mem_cp['o7101]='o0007;
mem_cp['o7102]='o7770;
mem_cp['o7103]='o0000;
mem_cp['o7104]='o0000;
mem_cp['o7105]='o0000;
mem_cp['o7106]='o0000;
mem_cp['o7107]='o0000;
mem_cp['o7110]='o0000;
mem_cp['o7111]='o0000;
mem_cp['o7112]='o0000;
mem_cp['o7113]='o0000;
mem_cp['o7114]='o0000;
mem_cp['o7115]='o0000;
mem_cp['o7116]='o0000;
mem_cp['o7117]='o0000;
mem_cp['o7120]='o0000;
mem_cp['o7121]='o0000;
mem_cp['o7122]='o0000;
mem_cp['o7123]='o0000;
mem_cp['o7124]='o0000;
mem_cp['o7125]='o0000;
mem_cp['o7126]='o0000;
mem_cp['o7127]='o0000;
mem_cp['o7130]='o0000;
mem_cp['o7131]='o0000;
mem_cp['o7132]='o0000;
mem_cp['o7133]='o0000;
mem_cp['o7134]='o0000;
mem_cp['o7135]='o0000;
mem_cp['o7136]='o0000;
mem_cp['o7137]='o0000;
mem_cp['o7140]='o0000;
mem_cp['o7141]='o0000;
mem_cp['o7142]='o0000;
mem_cp['o7143]='o0000;
mem_cp['o7144]='o0000;
mem_cp['o7145]='o0000;
mem_cp['o7146]='o0000;
mem_cp['o7147]='o0000;
mem_cp['o7150]='o0000;
mem_cp['o7151]='o0000;
mem_cp['o7152]='o0000;
mem_cp['o7153]='o0000;
mem_cp['o7154]='o0000;
mem_cp['o7155]='o0000;
mem_cp['o7156]='o0000;
mem_cp['o7157]='o0000;
mem_cp['o7160]='o0000;
mem_cp['o7161]='o0000;
mem_cp['o7162]='o0000;
mem_cp['o7163]='o0000;
mem_cp['o7164]='o0000;
mem_cp['o7165]='o0000;
mem_cp['o7166]='o0000;
mem_cp['o7167]='o0000;
mem_cp['o7170]='o0000;
mem_cp['o7171]='o0000;
mem_cp['o7172]='o0000;
mem_cp['o7173]='o0000;
mem_cp['o7174]='o0000;
mem_cp['o7175]='o0000;
mem_cp['o7176]='o0000;
mem_cp['o7177]='o0000;
mem_cp['o7200]='o0000;
mem_cp['o7201]='o7200;
mem_cp['o7202]='o1417;
mem_cp['o7203]='o7200;
mem_cp['o7204]='o1017;
mem_cp['o7205]='o0373;
mem_cp['o7206]='o1374;
mem_cp['o7207]='o3210;
mem_cp['o7210]='o7000;
mem_cp['o7211]='o7450;
mem_cp['o7212]='o5600;
mem_cp['o7213]='o3144;
mem_cp['o7214]='o4502;
mem_cp['o7215]='o5202;
mem_cp['o7216]='o0000;
mem_cp['o7217]='o7200;
mem_cp['o7220]='o1017;
mem_cp['o7221]='o3146;
mem_cp['o7222]='o4514;
mem_cp['o7223]='o4515;
mem_cp['o7224]='o5616;
mem_cp['o7225]='o0015;
mem_cp['o7226]='o0012;
mem_cp['o7227]='o0125;
mem_cp['o7230]='o0156;
mem_cp['o7231]='o0151;
mem_cp['o7232]='o0166;
mem_cp['o7233]='o0145;
mem_cp['o7234]='o0162;
mem_cp['o7235]='o0163;
mem_cp['o7236]='o0141;
mem_cp['o7237]='o0154;
mem_cp['o7240]='o0040;
mem_cp['o7241]='o0115;
mem_cp['o7242]='o0157;
mem_cp['o7243]='o0156;
mem_cp['o7244]='o0151;
mem_cp['o7245]='o0164;
mem_cp['o7246]='o0157;
mem_cp['o7247]='o0162;
mem_cp['o7250]='o0040;
mem_cp['o7251]='o0111;
mem_cp['o7252]='o0115;
mem_cp['o7253]='o0066;
mem_cp['o7254]='o0061;
mem_cp['o7255]='o0060;
mem_cp['o7256]='o0060;
mem_cp['o7257]='o0040;
mem_cp['o7260]='o0050;
mem_cp['o7261]='o0103;
mem_cp['o7262]='o0157;
mem_cp['o7263]='o0156;
mem_cp['o7264]='o0164;
mem_cp['o7265]='o0162;
mem_cp['o7266]='o0157;
mem_cp['o7267]='o0154;
mem_cp['o7270]='o0040;
mem_cp['o7271]='o0120;
mem_cp['o7272]='o0141;
mem_cp['o7273]='o0156;
mem_cp['o7274]='o0145;
mem_cp['o7275]='o0154;
mem_cp['o7276]='o0051;
mem_cp['o7277]='o0015;
mem_cp['o7300]='o0012;
mem_cp['o7301]='o0000;
mem_cp['o7302]='o0135;
mem_cp['o7303]='o0040;
mem_cp['o7304]='o0000;
mem_cp['o7305]='o0105;
mem_cp['o7306]='o0162;
mem_cp['o7307]='o0162;
mem_cp['o7310]='o0157;
mem_cp['o7311]='o0162;
mem_cp['o7312]='o0040;
mem_cp['o7313]='o0151;
mem_cp['o7314]='o0150;
mem_cp['o7315]='o0145;
mem_cp['o7316]='o0170;
mem_cp['o7317]='o0015;
mem_cp['o7320]='o0012;
mem_cp['o7321]='o0000;
mem_cp['o7322]='o0105;
mem_cp['o7323]='o0162;
mem_cp['o7324]='o0162;
mem_cp['o7325]='o0157;
mem_cp['o7326]='o0162;
mem_cp['o7327]='o0015;
mem_cp['o7330]='o0012;
mem_cp['o7331]='o0000;
mem_cp['o7332]='o0040;
mem_cp['o7333]='o0072;
mem_cp['o7334]='o0000;
mem_cp['o7335]='o0040;
mem_cp['o7336]='o0072;
mem_cp['o7337]='o0040;
mem_cp['o7340]='o0000;
mem_cp['o7341]='o0040;
mem_cp['o7342]='o0040;
mem_cp['o7343]='o0040;
mem_cp['o7344]='o0040;
mem_cp['o7345]='o0000;
mem_cp['o7346]='o0101;
mem_cp['o7347]='o0103;
mem_cp['o7350]='o0075;
mem_cp['o7351]='o0000;
mem_cp['o7352]='o0040;
mem_cp['o7353]='o0106;
mem_cp['o7354]='o0114;
mem_cp['o7355]='o0107;
mem_cp['o7356]='o0054;
mem_cp['o7357]='o0111;
mem_cp['o7360]='o0106;
mem_cp['o7361]='o0054;
mem_cp['o7362]='o0104;
mem_cp['o7363]='o0106;
mem_cp['o7364]='o0075;
mem_cp['o7365]='o0000;
mem_cp['o7366]='o0040;
mem_cp['o7367]='o0123;
mem_cp['o7370]='o0122;
mem_cp['o7371]='o0075;
mem_cp['o7372]='o0000;
mem_cp['o7373]='o0177;
mem_cp['o7374]='o1200;
mem_cp['o7375]='o0000;
mem_cp['o7376]='o0000;
mem_cp['o7377]='o0000;
mem_cp['o7400]='o0000;
mem_cp['o7401]='o6032;
mem_cp['o7402]='o6040;
mem_cp['o7403]='o7200;
mem_cp['o7404]='o5600;
mem_cp['o7405]='o0000;
mem_cp['o7406]='o6031;
mem_cp['o7407]='o5206;
mem_cp['o7410]='o6036;
mem_cp['o7411]='o0233;
mem_cp['o7412]='o3144;
mem_cp['o7413]='o5605;
mem_cp['o7414]='o0000;
mem_cp['o7415]='o7200;
mem_cp['o7416]='o7001;
mem_cp['o7417]='o6031;
mem_cp['o7420]='o7200;
mem_cp['o7421]='o3144;
mem_cp['o7422]='o5614;
mem_cp['o7423]='o0000;
mem_cp['o7424]='o6041;
mem_cp['o7425]='o5224;
mem_cp['o7426]='o7200;
mem_cp['o7427]='o1144;
mem_cp['o7430]='o6046;
mem_cp['o7431]='o7200;
mem_cp['o7432]='o5623;
mem_cp['o7433]='o0177;
mem_cp['o7434]='o0000;
mem_cp['o7435]='o0000;
mem_cp['o7436]='o0000;
mem_cp['o7437]='o0000;
mem_cp['o7440]='o0000;
mem_cp['o7441]='o0000;
mem_cp['o7442]='o0000;
mem_cp['o7443]='o0000;
mem_cp['o7444]='o0000;
mem_cp['o7445]='o0000;
mem_cp['o7446]='o0000;
mem_cp['o7447]='o0000;
mem_cp['o7450]='o0000;
mem_cp['o7451]='o0000;
mem_cp['o7452]='o0000;
mem_cp['o7453]='o0000;
mem_cp['o7454]='o0000;
mem_cp['o7455]='o0000;
mem_cp['o7456]='o0000;
mem_cp['o7457]='o0000;
mem_cp['o7460]='o0000;
mem_cp['o7461]='o0000;
mem_cp['o7462]='o0000;
mem_cp['o7463]='o0000;
mem_cp['o7464]='o0000;
mem_cp['o7465]='o0000;
mem_cp['o7466]='o0000;
mem_cp['o7467]='o0000;
mem_cp['o7470]='o0000;
mem_cp['o7471]='o0000;
mem_cp['o7472]='o0000;
mem_cp['o7473]='o0000;
mem_cp['o7474]='o0000;
mem_cp['o7475]='o0000;
mem_cp['o7476]='o0000;
mem_cp['o7477]='o0000;
mem_cp['o7500]='o0000;
mem_cp['o7501]='o0000;
mem_cp['o7502]='o0000;
mem_cp['o7503]='o0000;
mem_cp['o7504]='o0000;
mem_cp['o7505]='o0000;
mem_cp['o7506]='o0000;
mem_cp['o7507]='o0000;
mem_cp['o7510]='o0000;
mem_cp['o7511]='o0000;
mem_cp['o7512]='o0000;
mem_cp['o7513]='o0000;
mem_cp['o7514]='o0000;
mem_cp['o7515]='o0000;
mem_cp['o7516]='o0000;
mem_cp['o7517]='o0000;
mem_cp['o7520]='o0000;
mem_cp['o7521]='o0000;
mem_cp['o7522]='o0000;
mem_cp['o7523]='o0000;
mem_cp['o7524]='o0000;
mem_cp['o7525]='o0000;
mem_cp['o7526]='o0000;
mem_cp['o7527]='o0000;
mem_cp['o7530]='o0000;
mem_cp['o7531]='o0000;
mem_cp['o7532]='o0000;
mem_cp['o7533]='o0000;
mem_cp['o7534]='o0000;
mem_cp['o7535]='o0000;
mem_cp['o7536]='o0000;
mem_cp['o7537]='o0000;
mem_cp['o7540]='o0000;
mem_cp['o7541]='o0000;
mem_cp['o7542]='o0000;
mem_cp['o7543]='o0000;
mem_cp['o7544]='o0000;
mem_cp['o7545]='o0000;
mem_cp['o7546]='o0000;
mem_cp['o7547]='o0000;
mem_cp['o7550]='o0000;
mem_cp['o7551]='o0000;
mem_cp['o7552]='o0000;
mem_cp['o7553]='o0000;
mem_cp['o7554]='o0000;
mem_cp['o7555]='o0000;
mem_cp['o7556]='o0000;
mem_cp['o7557]='o0000;
mem_cp['o7560]='o0000;
mem_cp['o7561]='o0000;
mem_cp['o7562]='o0000;
mem_cp['o7563]='o0000;
mem_cp['o7564]='o0000;
mem_cp['o7565]='o0000;
mem_cp['o7566]='o0000;
mem_cp['o7567]='o0000;
mem_cp['o7570]='o0000;
mem_cp['o7571]='o0000;
mem_cp['o7572]='o0000;
mem_cp['o7573]='o0000;
mem_cp['o7574]='o0000;
mem_cp['o7575]='o0000;
mem_cp['o7576]='o0000;
mem_cp['o7577]='o0000;
mem_cp['o7600]='o0000;
mem_cp['o7601]='o0000;
mem_cp['o7602]='o0000;
mem_cp['o7603]='o0000;
mem_cp['o7604]='o0000;
mem_cp['o7605]='o0000;
mem_cp['o7606]='o0000;
mem_cp['o7607]='o0000;
mem_cp['o7610]='o0000;
mem_cp['o7611]='o0000;
mem_cp['o7612]='o0000;
mem_cp['o7613]='o0000;
mem_cp['o7614]='o0000;
mem_cp['o7615]='o0000;
mem_cp['o7616]='o0000;
mem_cp['o7617]='o0000;
mem_cp['o7620]='o0000;
mem_cp['o7621]='o0000;
mem_cp['o7622]='o0000;
mem_cp['o7623]='o0000;
mem_cp['o7624]='o0000;
mem_cp['o7625]='o0000;
mem_cp['o7626]='o0000;
mem_cp['o7627]='o0000;
mem_cp['o7630]='o0000;
mem_cp['o7631]='o0000;
mem_cp['o7632]='o0000;
mem_cp['o7633]='o0000;
mem_cp['o7634]='o0000;
mem_cp['o7635]='o0000;
mem_cp['o7636]='o0000;
mem_cp['o7637]='o0000;
mem_cp['o7640]='o0000;
mem_cp['o7641]='o0000;
mem_cp['o7642]='o0000;
mem_cp['o7643]='o0000;
mem_cp['o7644]='o0000;
mem_cp['o7645]='o0000;
mem_cp['o7646]='o0000;
mem_cp['o7647]='o0000;
mem_cp['o7650]='o0000;
mem_cp['o7651]='o0000;
mem_cp['o7652]='o0000;
mem_cp['o7653]='o0000;
mem_cp['o7654]='o0000;
mem_cp['o7655]='o0000;
mem_cp['o7656]='o0000;
mem_cp['o7657]='o0000;
mem_cp['o7660]='o0000;
mem_cp['o7661]='o0000;
mem_cp['o7662]='o0000;
mem_cp['o7663]='o0000;
mem_cp['o7664]='o0000;
mem_cp['o7665]='o0000;
mem_cp['o7666]='o0000;
mem_cp['o7667]='o0000;
mem_cp['o7670]='o0000;
mem_cp['o7671]='o0000;
mem_cp['o7672]='o0000;
mem_cp['o7673]='o0000;
mem_cp['o7674]='o0000;
mem_cp['o7675]='o0000;
mem_cp['o7676]='o0000;
mem_cp['o7677]='o0000;
mem_cp['o7700]='o0000;
mem_cp['o7701]='o0000;
mem_cp['o7702]='o0000;
mem_cp['o7703]='o0000;
mem_cp['o7704]='o0000;
mem_cp['o7705]='o0000;
mem_cp['o7706]='o0000;
mem_cp['o7707]='o0000;
mem_cp['o7710]='o0000;
mem_cp['o7711]='o0000;
mem_cp['o7712]='o0000;
mem_cp['o7713]='o0000;
mem_cp['o7714]='o0000;
mem_cp['o7715]='o0000;
mem_cp['o7716]='o0000;
mem_cp['o7717]='o0000;
mem_cp['o7720]='o0000;
mem_cp['o7721]='o0000;
mem_cp['o7722]='o0000;
mem_cp['o7723]='o0000;
mem_cp['o7724]='o0000;
mem_cp['o7725]='o0000;
mem_cp['o7726]='o0000;
mem_cp['o7727]='o0000;
mem_cp['o7730]='o0000;
mem_cp['o7731]='o0000;
mem_cp['o7732]='o0000;
mem_cp['o7733]='o0000;
mem_cp['o7734]='o0000;
mem_cp['o7735]='o0000;
mem_cp['o7736]='o0000;
mem_cp['o7737]='o0000;
mem_cp['o7740]='o0000;
mem_cp['o7741]='o0000;
mem_cp['o7742]='o0000;
mem_cp['o7743]='o0000;
mem_cp['o7744]='o0000;
mem_cp['o7745]='o0000;
mem_cp['o7746]='o0000;
mem_cp['o7747]='o0000;
mem_cp['o7750]='o0000;
mem_cp['o7751]='o0000;
mem_cp['o7752]='o0000;
mem_cp['o7753]='o0000;
mem_cp['o7754]='o0000;
mem_cp['o7755]='o0000;
mem_cp['o7756]='o0000;
mem_cp['o7757]='o0000;
mem_cp['o7760]='o0000;
mem_cp['o7761]='o0000;
mem_cp['o7762]='o0000;
mem_cp['o7763]='o0000;
mem_cp['o7764]='o0000;
mem_cp['o7765]='o0000;
mem_cp['o7766]='o0000;
mem_cp['o7767]='o0000;
mem_cp['o7770]='o0000;
mem_cp['o7771]='o0000;
mem_cp['o7772]='o0000;
mem_cp['o7773]='o0000;
mem_cp['o7774]='o0000;
mem_cp['o7775]='o0000;
mem_cp['o7776]='o5000;
mem_cp['o7777]='o5776;
end
